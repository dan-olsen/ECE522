
module dff_210 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_0 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_1 ( CK, Q, D );
  input CK, D;
  output Q;
  wire   n1;

  DFFX1 Q_reg ( .D(D), .CLK(CK), .QN(n1) );
  INVX0 U3 ( .INP(n1), .ZN(Q) );
endmodule


module dff_2 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_3 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_4 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_5 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_6 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_7 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_8 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_9 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_10 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_11 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_12 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_13 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_14 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_15 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_16 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_17 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_18 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_19 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_20 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_21 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_22 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_23 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_24 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_25 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_26 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_27 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_28 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_29 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_30 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_31 ( CK, Q, D );
  input CK, D;
  output Q;
  wire   n1;

  DFFX2 Q_reg ( .D(D), .CLK(CK), .QN(n1) );
  INVX0 U3 ( .INP(n1), .ZN(Q) );
endmodule


module dff_32 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_33 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_34 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_35 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_36 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_37 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_38 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_39 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_40 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_41 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_42 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_43 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_44 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_45 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_46 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_47 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_48 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_49 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_50 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_51 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_52 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_53 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_54 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_55 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_56 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_57 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_58 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_59 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_60 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_61 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_62 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_63 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_64 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_65 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_66 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_67 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_68 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_69 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_70 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_71 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_72 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_73 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_74 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_75 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_76 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_77 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_78 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_79 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_80 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_81 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_82 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_83 ( CK, Q, D );
  input CK, D;
  output Q;
  wire   n1;

  DFFX1 Q_reg ( .D(D), .CLK(CK), .QN(n1) );
  INVX0 U3 ( .INP(n1), .ZN(Q) );
endmodule


module dff_84 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_85 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_86 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_87 ( CK, Q, D );
  input CK, D;
  output Q;
  wire   n1;

  DFFX2 Q_reg ( .D(D), .CLK(CK), .QN(n1) );
  INVX1 U3 ( .INP(n1), .ZN(Q) );
endmodule


module dff_88 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_89 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_90 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_91 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_92 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_93 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_94 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_95 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_96 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_97 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_98 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_99 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_100 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_101 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_102 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_103 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_104 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_105 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_106 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_107 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_108 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_109 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_110 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_111 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_112 ( CK, Q, D );
  input CK, D;
  output Q;
  wire   n1;

  DFFX2 Q_reg ( .D(D), .CLK(CK), .QN(n1) );
  INVX0 U3 ( .INP(n1), .ZN(Q) );
endmodule


module dff_113 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_114 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_115 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_116 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_117 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_118 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_119 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_120 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_121 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_122 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_123 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_124 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_125 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_126 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_127 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_128 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_129 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_130 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_131 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_132 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_133 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_134 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_135 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_136 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_137 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_138 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_139 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_140 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_141 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_142 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_143 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_144 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_145 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_146 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_147 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_148 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_149 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_150 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_151 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_152 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_153 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_154 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_155 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_156 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_157 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_158 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_159 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_160 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_161 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_162 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_163 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_164 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_165 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_166 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_167 ( CK, Q, D );
  input CK, D;
  output Q;
  wire   n1;

  DFFX2 Q_reg ( .D(D), .CLK(CK), .QN(n1) );
  INVX0 U3 ( .INP(n1), .ZN(Q) );
endmodule


module dff_168 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_169 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_170 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_171 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_172 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_173 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_174 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_175 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_176 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_177 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_178 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_179 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_180 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_181 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_182 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_183 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_184 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_185 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_186 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_187 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_188 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_189 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_190 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_191 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_192 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_193 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_194 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_195 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_196 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_197 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_198 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_199 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_200 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_201 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_202 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_203 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_204 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_205 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_206 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_207 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_208 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module dff_209 ( CK, Q, D );
  input CK, D;
  output Q;


  DFFX1 Q_reg ( .D(D), .CLK(CK), .Q(Q) );
endmodule


module s9234 ( CK, g102, g107, g1290, g1293, g22, g23, g2584, g301, g306, g310, 
        g314, g319, g32, g3222, g36, g3600, g37, g38, g39, g40, g4098, g4099, 
        g41, g4100, g4101, g4102, g4103, g4104, g4105, g4106, g4107, g4108, 
        g4109, g4110, g4112, g4121, g42, g4307, g4321, g44, g4422, g45, g46, 
        g47, g4809, g5137, g5468, g5469, g557, g558, g559, g560, g561, g562, 
        g563, g564, g567, g5692, g6282, g6284, g6360, g6362, g6364, g6366, 
        g6368, g6370, g6372, g6374, g639, g6728, g702, g705, g89, g94, g98 );
  input CK, g102, g107, g22, g23, g301, g306, g310, g314, g319, g32, g36, g37,
         g38, g39, g40, g41, g42, g44, g45, g46, g47, g557, g558, g559, g560,
         g561, g562, g563, g564, g567, g639, g702, g705, g89, g94, g98;
  output g1290, g1293, g2584, g3222, g3600, g4098, g4099, g4100, g4101, g4102,
         g4103, g4104, g4105, g4106, g4107, g4108, g4109, g4110, g4112, g4121,
         g4307, g4321, g4422, g4809, g5137, g5468, g5469, g5692, g6282, g6284,
         g6360, g6362, g6364, g6366, g6368, g6370, g6372, g6374, g6728;
  wire   g678, g332, g123, g207, g695, g461, g18, g292, g331, g689, g24, g465,
         g84, g291, g676, g622, g117, g278, g128, g598, g554, g496, g179, g48,
         g590, g551, g682, g606, g188, g646, g327, g361, g289, g398, g5700,
         g684, g619, g208, g248, g390, g5698, g625, g681, g437, g276, g323,
         g224, g685, g43, g157, g5470, g282, g697, g206, g449, g118, g528,
         g284, g426, g634, g669, g520, g281, g175, g5472, g631, g69, g693,
         g337, g457, g486, g471, g328, g285, g418, g402, g297, g212, g410,
         g430, g662, g453, g269, g574, g441, g664, g349, g211, g586, g571,
         g326, g698, g654, g293, g690, g445, g374, g5694, g6, g687, g357, g386,
         g5697, g504, g665, g166, g5471, g541, g74, g338, g696, g516, g536,
         g683, g353, g545, g254, g341, g290, g2, g287, g336, g345, g628, g679,
         g28, g688, g283, g613, g10, g14, g680, g143, g672, g667, g366, g279,
         g492, g170, g686, g288, g638, g602, g642, g280, g663, g610, g148,
         g209, g675, g478, g122, g54, g594, g286, g489, g616, g79, g218, g242,
         g578, g184, g5473, g119, g668, g139, g422, g210, g394, g5699, g230,
         g204, g658, g650, g378, g5695, g508, g548, g370, g5693, g406, g236,
         g500, g205, g197, g666, g114, g524, g260, g111, g131, g677, g582,
         g485, g699, g193, g5474, g135, g382, g5696, g414, g434, g266, g49,
         g152, g692, g277, g127, g161, g512, g532, g64, g694, g691, g1, g59,
         g5624, g6294, g5386, g6688, g6110, g6300, g6485, g4757, g6173, g6182,
         g6426, g4430, g2859, g6795, g6686, g3725, g4446, g6292, g6689, g6481,
         g6297, g5231, g5531, g3729, g5626, g4447, g3731, g2670, g6293, g6690,
         g6179, g6791, g6691, g6794, g6453, g6113, g6167, g4444, g5627, g6792,
         g6286, g5630, g6684, g4740, g6109, g4458, g6307, g4454, g5916, g6658,
         g5628, g3727, g6455, g5291, g4433, g6845, g6483, g4219, g6176, g3724,
         g6299, g6142, g6704, g4752, g6309, g6787, g6454, g6456, g4872, g4497,
         g6296, g5625, g4460, g3768, g6793, g4607, g4501, g4440, g6790, g6452,
         g6185, g4436, g3828, g6310, g6687, g5629, g6937, g3454, g6921, g6301,
         g5532, g4441, g4157, g3730, g5303, g5533, g6170, g5277, g4443, g6304,
         g6844, g6189, g6116, g5583, g4761, g5535, g5622, g6480, g6447, g6298,
         g2433, g6290, g6114, g4451, g6685, g6450, g6437, g6789, g6291, g5323,
         g3728, g6444, g5295, g6118, g2861, g5050, g4434, g4687, g6108, g6287,
         g3844, g4438, g1802, g3726, g6482, g5017, g3910, g6303, g6440, g5149,
         g5701, g6788, g6702, g4773, g6936, g4450, g3814, g6295, g5167, g4455,
         g3599, g6289, g6479, n2, n3, n4, n6, n8, n11, n12, n13, n14, n15, n16,
         n17, n18, n20, n21, n23, n24, n26, n27, n28, n29, n31, n32, n33, n34,
         n35, n37, n38, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n66, n67,
         n68, n69, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n94, n95, n96, n97,
         n99, n100, n101, n102, n103, n104, n105, n106, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n143, n144, n145,
         n147, n148, n151, n152, n154, n155, n156, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n255, n256, n260, n261, n263, n264, n265, n266, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n288, n291, n292, n293, n294, n295, n296,
         n297, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n361, n362, n363, n364, n366, n367,
         n368, n369, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n406, n407, n408, n409, n410, n412, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n508, n509, n511,
         n512, n513, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n536, n537,
         n538, n539, n540, n541, n542, n543, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n582, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n603, n604, n605, n606, n607, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n726, n728, n730,
         n732, n734, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n938, n940, n942, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046;
  assign g3600 = g43;
  assign g4321 = g668;
  assign g1290 = g666;
  assign g4307 = g485;
  assign g6284 = g6110;
  assign g6370 = g6173;
  assign g6360 = g6182;
  assign g6374 = g6179;
  assign g6364 = g6167;
  assign g6372 = g6176;
  assign g6362 = g6185;
  assign g6368 = g6170;
  assign g6366 = g6189;
  assign g4809 = g2433;
  assign g2584 = g1802;
  assign g4121 = g3599;

  dff_210 DFF_0 ( .CK(CK), .Q(g678), .D(n824) );
  dff_209 DFF_1 ( .CK(CK), .Q(g332), .D(g6795) );
  dff_208 DFF_2 ( .CK(CK), .Q(g123), .D(g6937) );
  dff_207 DFF_3 ( .CK(CK), .Q(g207), .D(g5626) );
  dff_206 DFF_4 ( .CK(CK), .Q(g695), .D(n812) );
  dff_205 DFF_5 ( .CK(CK), .Q(g461), .D(g4440) );
  dff_204 DFF_6 ( .CK(CK), .Q(g18), .D(g6684) );
  dff_203 DFF_7 ( .CK(CK), .Q(g292), .D(g571) );
  dff_202 DFF_8 ( .CK(CK), .Q(g331), .D(g3730) );
  dff_201 DFF_9 ( .CK(CK), .Q(g689), .D(g4103) );
  dff_200 DFF_10 ( .CK(CK), .Q(g24), .D(g6685) );
  dff_199 DFF_11 ( .CK(CK), .Q(g465), .D(g6297) );
  dff_198 DFF_12 ( .CK(CK), .Q(g84), .D(g6456) );
  dff_197 DFF_13 ( .CK(CK), .Q(g291), .D(g654) );
  dff_196 DFF_14 ( .CK(CK), .Q(g676), .D(n23) );
  dff_195 DFF_15 ( .CK(CK), .Q(g622), .D(g4460) );
  dff_194 DFF_16 ( .CK(CK), .Q(g117), .D(g4497) );
  dff_193 DFF_17 ( .CK(CK), .Q(g278), .D(g5627) );
  dff_192 DFF_18 ( .CK(CK), .Q(g128), .D(g4773) );
  dff_191 DFF_19 ( .CK(CK), .Q(g598), .D(g2859) );
  dff_190 DFF_20 ( .CK(CK), .Q(g554), .D(g6790) );
  dff_189 DFF_21 ( .CK(CK), .Q(g496), .D(g6702) );
  dff_188 DFF_22 ( .CK(CK), .Q(g179), .D(g6116) );
  dff_187 DFF_23 ( .CK(CK), .Q(g48), .D(g6658) );
  dff_186 DFF_24 ( .CK(CK), .Q(g590), .D(g6437) );
  dff_185 DFF_25 ( .CK(CK), .Q(g551), .D(g6789) );
  dff_184 DFF_26 ( .CK(CK), .Q(g682), .D(n812) );
  dff_183 DFF_27 ( .CK(CK), .Q(g6689), .D(g6481) );
  dff_182 DFF_28 ( .CK(CK), .Q(g606), .D(g4219) );
  dff_181 DFF_29 ( .CK(CK), .Q(g188), .D(g6118) );
  dff_180 DFF_30 ( .CK(CK), .Q(g646), .D(g4501) );
  dff_179 DFF_31 ( .CK(CK), .Q(g327), .D(g3728) );
  dff_178 DFF_32 ( .CK(CK), .Q(g361), .D(g6440) );
  dff_177 DFF_33 ( .CK(CK), .Q(g289), .D(g646) );
  dff_176 DFF_34 ( .CK(CK), .Q(g398), .D(g5700) );
  dff_175 DFF_35 ( .CK(CK), .Q(g684), .D(n825) );
  dff_174 DFF_36 ( .CK(CK), .Q(g619), .D(g4157) );
  dff_173 DFF_37 ( .CK(CK), .Q(g208), .D(g5533) );
  dff_172 DFF_38 ( .CK(CK), .Q(g248), .D(g650) );
  dff_171 DFF_39 ( .CK(CK), .Q(g390), .D(g5698) );
  dff_170 DFF_40 ( .CK(CK), .Q(g625), .D(g4687) );
  dff_169 DFF_41 ( .CK(CK), .Q(g681), .D(n815) );
  dff_168 DFF_42 ( .CK(CK), .Q(g437), .D(g4433) );
  dff_167 DFF_43 ( .CK(CK), .Q(g276), .D(g5532) );
  dff_166 DFF_44 ( .CK(CK), .Q(g6686), .D(g6479) );
  dff_165 DFF_45 ( .CK(CK), .Q(g323), .D(g3731) );
  dff_164 DFF_46 ( .CK(CK), .Q(g224), .D(n892) );
  dff_163 DFF_47 ( .CK(CK), .Q(g685), .D(g4099) );
  dff_162 DFF_48 ( .CK(CK), .Q(g43), .D(g6142) );
  dff_161 DFF_49 ( .CK(CK), .Q(g157), .D(g5470) );
  dff_160 DFF_50 ( .CK(CK), .Q(g282), .D(g6793) );
  dff_159 DFF_51 ( .CK(CK), .Q(g697), .D(n825) );
  dff_158 DFF_52 ( .CK(CK), .Q(g206), .D(g5624) );
  dff_157 DFF_53 ( .CK(CK), .Q(g449), .D(g4450) );
  dff_156 DFF_54 ( .CK(CK), .Q(g118), .D(g3724) );
  dff_155 DFF_55 ( .CK(CK), .Q(g528), .D(g6286) );
  dff_154 DFF_56 ( .CK(CK), .Q(g284), .D(n986) );
  dff_153 DFF_57 ( .CK(CK), .Q(g426), .D(g4458) );
  dff_152 DFF_58 ( .CK(CK), .Q(g634), .D(g3454) );
  dff_151 DFF_59 ( .CK(CK), .Q(g669), .D(g5386) );
  dff_150 DFF_60 ( .CK(CK), .Q(g520), .D(g6309) );
  dff_149 DFF_61 ( .CK(CK), .Q(g281), .D(g5630) );
  dff_148 DFF_62 ( .CK(CK), .Q(g175), .D(g5472) );
  dff_147 DFF_63 ( .CK(CK), .Q(g6690), .D(g6482) );
  dff_146 DFF_64 ( .CK(CK), .Q(g631), .D(g5167) );
  dff_145 DFF_65 ( .CK(CK), .Q(g69), .D(g6453) );
  dff_144 DFF_66 ( .CK(CK), .Q(g693), .D(n816) );
  dff_143 DFF_67 ( .CK(CK), .Q(g337), .D(n148) );
  dff_142 DFF_68 ( .CK(CK), .Q(g457), .D(g4443) );
  dff_141 DFF_69 ( .CK(CK), .Q(g486), .D(n980) );
  dff_140 DFF_70 ( .CK(CK), .Q(g471), .D(g664) );
  dff_139 DFF_71 ( .CK(CK), .Q(g328), .D(g3729) );
  dff_138 DFF_72 ( .CK(CK), .Q(g285), .D(n966) );
  dff_137 DFF_73 ( .CK(CK), .Q(g418), .D(g4451) );
  dff_136 DFF_74 ( .CK(CK), .Q(g402), .D(g4438) );
  dff_135 DFF_75 ( .CK(CK), .Q(g297), .D(g6298) );
  dff_134 DFF_76 ( .CK(CK), .Q(g212), .D(n985) );
  dff_133 DFF_77 ( .CK(CK), .Q(g410), .D(g4444) );
  dff_132 DFF_78 ( .CK(CK), .Q(g430), .D(g4434) );
  dff_131 DFF_79 ( .CK(CK), .Q(g6687), .D(g6845) );
  dff_130 DFF_80 ( .CK(CK), .Q(g662), .D(n131) );
  dff_129 DFF_81 ( .CK(CK), .Q(g453), .D(g4446) );
  dff_128 DFF_82 ( .CK(CK), .Q(g269), .D(g6290) );
  dff_127 DFF_83 ( .CK(CK), .Q(g574), .D(g6426) );
  dff_126 DFF_84 ( .CK(CK), .Q(g441), .D(g4430) );
  dff_125 DFF_85 ( .CK(CK), .Q(g664), .D(g663) );
  dff_124 DFF_86 ( .CK(CK), .Q(g349), .D(g5295) );
  dff_123 DFF_87 ( .CK(CK), .Q(g211), .D(g6792) );
  dff_122 DFF_88 ( .CK(CK), .Q(g586), .D(g6299) );
  dff_121 DFF_89 ( .CK(CK), .Q(g571), .D(g5149) );
  dff_120 DFF_90 ( .CK(CK), .Q(g6685), .D(g6844) );
  dff_119 DFF_91 ( .CK(CK), .Q(g326), .D(g4607) );
  dff_118 DFF_92 ( .CK(CK), .Q(g698), .D(g4105) );
  dff_117 DFF_93 ( .CK(CK), .Q(g654), .D(g5017) );
  dff_116 DFF_94 ( .CK(CK), .Q(g293), .D(g6294) );
  dff_115 DFF_95 ( .CK(CK), .Q(g690), .D(n817) );
  dff_114 DFF_96 ( .CK(CK), .Q(g445), .D(g4454) );
  dff_113 DFF_97 ( .CK(CK), .Q(g374), .D(g5694) );
  dff_112 DFF_98 ( .CK(CK), .Q(g6), .D(g6689) );
  dff_111 DFF_99 ( .CK(CK), .Q(g687), .D(g4101) );
  dff_110 DFF_100 ( .CK(CK), .Q(g357), .D(g5303) );
  dff_109 DFF_101 ( .CK(CK), .Q(g386), .D(g5697) );
  dff_108 DFF_102 ( .CK(CK), .Q(g504), .D(g6296) );
  dff_107 DFF_103 ( .CK(CK), .Q(g665), .D(g42) );
  dff_106 DFF_104 ( .CK(CK), .Q(g166), .D(g5471) );
  dff_105 DFF_105 ( .CK(CK), .Q(g541), .D(g6289) );
  dff_104 DFF_106 ( .CK(CK), .Q(g74), .D(g6454) );
  dff_103 DFF_107 ( .CK(CK), .Q(g338), .D(g5323) );
  dff_102 DFF_108 ( .CK(CK), .Q(g696), .D(n818) );
  dff_101 DFF_109 ( .CK(CK), .Q(g516), .D(g6307) );
  dff_100 DFF_110 ( .CK(CK), .Q(g536), .D(g6293) );
  dff_99 DFF_111 ( .CK(CK), .Q(g683), .D(n818) );
  dff_98 DFF_112 ( .CK(CK), .Q(g353), .D(g5050) );
  dff_97 DFF_113 ( .CK(CK), .Q(g545), .D(g6787) );
  dff_96 DFF_114 ( .CK(CK), .Q(g254), .D(g654) );
  dff_95 DFF_115 ( .CK(CK), .Q(g341), .D(g5277) );
  dff_94 DFF_116 ( .CK(CK), .Q(g290), .D(g650) );
  dff_93 DFF_117 ( .CK(CK), .Q(g2), .D(g6688) );
  dff_92 DFF_118 ( .CK(CK), .Q(g287), .D(n720) );
  dff_91 DFF_119 ( .CK(CK), .Q(g336), .D(g6921) );
  dff_90 DFF_120 ( .CK(CK), .Q(g345), .D(g5291) );
  dff_89 DFF_121 ( .CK(CK), .Q(g628), .D(g4872) );
  dff_88 DFF_122 ( .CK(CK), .Q(g679), .D(n823) );
  dff_87 DFF_123 ( .CK(CK), .Q(g28), .D(g6687) );
  dff_86 DFF_124 ( .CK(CK), .Q(g688), .D(g4102) );
  dff_85 DFF_125 ( .CK(CK), .Q(g283), .D(n1019) );
  dff_84 DFF_126 ( .CK(CK), .Q(g613), .D(g3828) );
  dff_83 DFF_127 ( .CK(CK), .Q(g10), .D(g6690) );
  dff_82 DFF_128 ( .CK(CK), .Q(g14), .D(g6691) );
  dff_81 DFF_129 ( .CK(CK), .Q(g680), .D(n816) );
  dff_80 DFF_130 ( .CK(CK), .Q(g143), .D(g6108) );
  dff_79 DFF_131 ( .CK(CK), .Q(g672), .D(g5231) );
  dff_78 DFF_132 ( .CK(CK), .Q(g667), .D(g45) );
  dff_77 DFF_133 ( .CK(CK), .Q(g366), .D(g5916) );
  dff_76 DFF_134 ( .CK(CK), .Q(g279), .D(g5628) );
  dff_75 DFF_135 ( .CK(CK), .Q(g492), .D(g6704) );
  dff_74 DFF_136 ( .CK(CK), .Q(g170), .D(g6114) );
  dff_73 DFF_137 ( .CK(CK), .Q(g686), .D(g4100) );
  dff_72 DFF_138 ( .CK(CK), .Q(g288), .D(n702) );
  dff_71 DFF_139 ( .CK(CK), .Q(g638), .D(g667) );
  dff_70 DFF_140 ( .CK(CK), .Q(g602), .D(g2861) );
  dff_69 DFF_141 ( .CK(CK), .Q(g642), .D(g3844) );
  dff_68 DFF_142 ( .CK(CK), .Q(g280), .D(g5535) );
  dff_67 DFF_143 ( .CK(CK), .Q(g663), .D(g42) );
  dff_66 DFF_144 ( .CK(CK), .Q(g610), .D(g2670) );
  dff_65 DFF_145 ( .CK(CK), .Q(g148), .D(g5583) );
  dff_64 DFF_146 ( .CK(CK), .Q(g209), .D(g5629) );
  dff_63 DFF_147 ( .CK(CK), .Q(g675), .D(g702) );
  dff_62 DFF_148 ( .CK(CK), .Q(g478), .D(g665) );
  dff_61 DFF_149 ( .CK(CK), .Q(g122), .D(g3726) );
  dff_60 DFF_150 ( .CK(CK), .Q(g54), .D(g6447) );
  dff_59 DFF_151 ( .CK(CK), .Q(g594), .D(g6304) );
  dff_58 DFF_152 ( .CK(CK), .Q(g286), .D(n892) );
  dff_57 DFF_153 ( .CK(CK), .Q(g489), .D(n136) );
  dff_56 DFF_154 ( .CK(CK), .Q(g616), .D(g3768) );
  dff_55 DFF_155 ( .CK(CK), .Q(g79), .D(g6455) );
  dff_54 DFF_156 ( .CK(CK), .Q(g218), .D(n965) );
  dff_53 DFF_157 ( .CK(CK), .Q(g242), .D(g646) );
  dff_52 DFF_158 ( .CK(CK), .Q(g578), .D(g6291) );
  dff_51 DFF_159 ( .CK(CK), .Q(g184), .D(g5473) );
  dff_50 DFF_160 ( .CK(CK), .Q(g119), .D(g3725) );
  dff_49 DFF_161 ( .CK(CK), .Q(g668), .D(n655) );
  dff_48 DFF_162 ( .CK(CK), .Q(g139), .D(g4757) );
  dff_47 DFF_163 ( .CK(CK), .Q(g422), .D(g4455) );
  dff_46 DFF_164 ( .CK(CK), .Q(g210), .D(g6791) );
  dff_45 DFF_165 ( .CK(CK), .Q(g394), .D(g5699) );
  dff_44 DFF_166 ( .CK(CK), .Q(g230), .D(n720) );
  dff_43 DFF_167 ( .CK(CK), .Q(g6684), .D(g6485) );
  dff_42 DFF_168 ( .CK(CK), .Q(g204), .D(g5531) );
  dff_41 DFF_169 ( .CK(CK), .Q(g658), .D(g3814) );
  dff_40 DFF_170 ( .CK(CK), .Q(g650), .D(g4761) );
  dff_39 DFF_171 ( .CK(CK), .Q(g378), .D(g5695) );
  dff_38 DFF_172 ( .CK(CK), .Q(g508), .D(g6300) );
  dff_37 DFF_173 ( .CK(CK), .Q(g548), .D(g6788) );
  dff_36 DFF_174 ( .CK(CK), .Q(g370), .D(g5693) );
  dff_35 DFF_175 ( .CK(CK), .Q(g406), .D(g4441) );
  dff_34 DFF_176 ( .CK(CK), .Q(g236), .D(n702) );
  dff_33 DFF_177 ( .CK(CK), .Q(g500), .D(g6292) );
  dff_32 DFF_178 ( .CK(CK), .Q(g205), .D(g5622) );
  dff_31 DFF_179 ( .CK(CK), .Q(g197), .D(g6287) );
  dff_30 DFF_180 ( .CK(CK), .Q(g666), .D(g46) );
  dff_29 DFF_181 ( .CK(CK), .Q(g114), .D(g3727) );
  dff_28 DFF_182 ( .CK(CK), .Q(g524), .D(g6310) );
  dff_27 DFF_183 ( .CK(CK), .Q(g260), .D(g571) );
  dff_26 DFF_184 ( .CK(CK), .Q(g111), .D(g5701) );
  dff_25 DFF_185 ( .CK(CK), .Q(g131), .D(g4740) );
  dff_24 DFF_186 ( .CK(CK), .Q(g6688), .D(g6480) );
  dff_23 DFF_187 ( .CK(CK), .Q(g6691), .D(g6483) );
  dff_22 DFF_188 ( .CK(CK), .Q(g677), .D(n817) );
  dff_21 DFF_189 ( .CK(CK), .Q(g582), .D(g6295) );
  dff_20 DFF_190 ( .CK(CK), .Q(g485), .D(n656) );
  dff_19 DFF_191 ( .CK(CK), .Q(g699), .D(n940) );
  dff_18 DFF_192 ( .CK(CK), .Q(g193), .D(g5474) );
  dff_17 DFF_193 ( .CK(CK), .Q(g135), .D(g4752) );
  dff_16 DFF_194 ( .CK(CK), .Q(g382), .D(g5696) );
  dff_15 DFF_195 ( .CK(CK), .Q(g414), .D(g4447) );
  dff_14 DFF_196 ( .CK(CK), .Q(g434), .D(g4436) );
  dff_13 DFF_197 ( .CK(CK), .Q(g266), .D(g3910) );
  dff_12 DFF_198 ( .CK(CK), .Q(g49), .D(g6444) );
  dff_11 DFF_199 ( .CK(CK), .Q(g152), .D(g6109) );
  dff_10 DFF_200 ( .CK(CK), .Q(g692), .D(n823) );
  dff_9 DFF_201 ( .CK(CK), .Q(g277), .D(g5625) );
  dff_8 DFF_202 ( .CK(CK), .Q(g127), .D(g6936) );
  dff_7 DFF_203 ( .CK(CK), .Q(g161), .D(g6113) );
  dff_6 DFF_204 ( .CK(CK), .Q(g512), .D(g6303) );
  dff_5 DFF_205 ( .CK(CK), .Q(g532), .D(g6301) );
  dff_4 DFF_206 ( .CK(CK), .Q(g64), .D(g6452) );
  dff_3 DFF_207 ( .CK(CK), .Q(g694), .D(n815) );
  dff_2 DFF_208 ( .CK(CK), .Q(g691), .D(n824) );
  dff_1 DFF_209 ( .CK(CK), .Q(g1), .D(g6686) );
  dff_0 DFF_210 ( .CK(CK), .Q(g59), .D(g6450) );
  NAND3X0 U341 ( .IN1(n168), .IN2(n169), .IN3(n170), .QN(n163) );
  AO221X1 U344 ( .IN1(n176), .IN2(g297), .IN3(n862), .IN4(n656), .IN5(n177), 
        .Q(n168) );
  AO22X1 U345 ( .IN1(n140), .IN2(n180), .IN3(n181), .IN4(n827), .Q(g6936) );
  AO22X1 U346 ( .IN1(n139), .IN2(n125), .IN3(g127), .IN4(n183), .Q(n181) );
  NAND4X0 U347 ( .IN1(n184), .IN2(g119), .IN3(n185), .IN4(n186), .QN(n183) );
  NAND4X0 U348 ( .IN1(n187), .IN2(n188), .IN3(n189), .IN4(n190), .QN(n185) );
  OA22X1 U350 ( .IN1(g123), .IN2(n187), .IN3(n11), .IN4(n190), .Q(n191) );
  AO221X1 U354 ( .IN1(n199), .IN2(n63), .IN3(n52), .IN4(n710), .IN5(n110), .Q(
        n197) );
  OAI221X1 U355 ( .IN1(n201), .IN2(g650), .IN3(n200), .IN4(g606), .IN5(g260), 
        .QN(n196) );
  AO22X1 U356 ( .IN1(g680), .IN2(n983), .IN3(g646), .IN4(n862), .Q(n200) );
  AO221X1 U361 ( .IN1(n176), .IN2(g293), .IN3(n967), .IN4(n655), .IN5(n177), 
        .Q(n194) );
  AO22X1 U362 ( .IN1(n981), .IN2(n983), .IN3(n204), .IN4(n968), .Q(n177) );
  OA22X1 U363 ( .IN1(n205), .IN2(n206), .IN3(n207), .IN4(n208), .Q(n204) );
  NAND4X0 U364 ( .IN1(n209), .IN2(n210), .IN3(n211), .IN4(n212), .QN(n208) );
  NAND4X0 U366 ( .IN1(n739), .IN2(n892), .IN3(n986), .IN4(n42), .QN(n211) );
  NAND4X0 U367 ( .IN1(g696), .IN2(n892), .IN3(n966), .IN4(n158), .QN(n210) );
  NAND4X0 U368 ( .IN1(n215), .IN2(n216), .IN3(n217), .IN4(n218), .QN(n207) );
  NAND3X0 U369 ( .IN1(g690), .IN2(n76), .IN3(n213), .QN(n218) );
  NAND4X0 U370 ( .IN1(g567), .IN2(g691), .IN3(n42), .IN4(n76), .QN(n217) );
  NAND4X0 U371 ( .IN1(n965), .IN2(g692), .IN3(n158), .IN4(n76), .QN(n216) );
  NAND4X0 U373 ( .IN1(n220), .IN2(n221), .IN3(n222), .IN4(n223), .QN(n206) );
  XOR2X1 U374 ( .IN1(n63), .IN2(g287), .Q(n223) );
  XNOR2X1 U375 ( .IN1(g680), .IN2(g286), .Q(n222) );
  XOR2X1 U376 ( .IN1(n710), .IN2(g285), .Q(n221) );
  XOR2X1 U377 ( .IN1(n4), .IN2(g284), .Q(n220) );
  NAND4X0 U378 ( .IN1(n224), .IN2(n225), .IN3(n226), .IN4(n227), .QN(n205) );
  XOR2X1 U380 ( .IN1(g686), .IN2(g292), .Q(n229) );
  XOR2X1 U382 ( .IN1(n100), .IN2(g289), .Q(n225) );
  XOR2X1 U383 ( .IN1(n48), .IN2(g288), .Q(n224) );
  AOI22X1 U384 ( .IN1(g254), .IN2(g248), .IN3(g242), .IN4(g236), .QN(n232) );
  AO22X1 U385 ( .IN1(n749), .IN2(n233), .IN3(n234), .IN4(n235), .Q(g6921) );
  AO21X1 U386 ( .IN1(g336), .IN2(n236), .IN3(n151), .Q(n234) );
  NAND4X0 U388 ( .IN1(n240), .IN2(n241), .IN3(n811), .IN4(n242), .QN(n238) );
  AND2X1 U391 ( .IN1(n703), .IN2(n244), .Q(n240) );
  NAND4X0 U392 ( .IN1(n247), .IN2(n246), .IN3(n245), .IN4(n248), .QN(n233) );
  AO221X1 U412 ( .IN1(n277), .IN2(n275), .IN3(n276), .IN4(n278), .IN5(n1017), 
        .Q(n273) );
  AO221X1 U415 ( .IN1(n281), .IN2(g683), .IN3(g685), .IN4(n282), .IN5(n992), 
        .Q(n246) );
  AO221X1 U416 ( .IN1(n277), .IN2(n281), .IN3(n282), .IN4(n278), .IN5(n1011), 
        .Q(n245) );
  AO22X1 U420 ( .IN1(g646), .IN2(n862), .IN3(g242), .IN4(n983), .Q(n277) );
  AO22X1 U422 ( .IN1(n702), .IN2(n968), .IN3(g236), .IN4(n983), .Q(n280) );
  AOI221X1 U424 ( .IN1(g6792), .IN2(n876), .IN3(n1019), .IN4(n679), .IN5(n288), 
        .QN(n286) );
  NAND4X0 U427 ( .IN1(n292), .IN2(n910), .IN3(n293), .IN4(n294), .QN(g6844) );
  AOI221X1 U428 ( .IN1(g6791), .IN2(n974), .IN3(g6793), .IN4(n979), .IN5(n295), 
        .QN(n294) );
  AO221X1 U438 ( .IN1(n302), .IN2(n857), .IN3(n303), .IN4(g283), .IN5(n16), 
        .Q(n179) );
  AOI21X1 U442 ( .IN1(n33), .IN2(g283), .IN3(n312), .QN(n303) );
  AO221X1 U444 ( .IN1(n313), .IN2(n852), .IN3(n314), .IN4(g211), .IN5(n15), 
        .Q(n231) );
  NAND3X0 U446 ( .IN1(n315), .IN2(n318), .IN3(g210), .QN(n317) );
  AND3X1 U447 ( .IN1(n321), .IN2(g210), .IN3(n322), .Q(n316) );
  AOI21X1 U448 ( .IN1(n14), .IN2(g211), .IN3(n323), .QN(n314) );
  NAND3X0 U449 ( .IN1(g282), .IN2(n325), .IN3(g283), .QN(n324) );
  AO22X1 U450 ( .IN1(n310), .IN2(n311), .IN3(n308), .IN4(n78), .Q(n325) );
  XOR2X1 U451 ( .IN1(g478), .IN2(n844), .Q(n308) );
  NAND4X0 U453 ( .IN1(g278), .IN2(n330), .IN3(n331), .IN4(n332), .QN(n329) );
  OR2X1 U455 ( .IN1(n917), .IN2(g690), .Q(n331) );
  AO221X1 U456 ( .IN1(g693), .IN2(n64), .IN3(n762), .IN4(g692), .IN5(n803), 
        .Q(n330) );
  OA22X1 U458 ( .IN1(n803), .IN2(n336), .IN3(g694), .IN4(n917), .Q(n335) );
  NAND3X0 U461 ( .IN1(g210), .IN2(n338), .IN3(g211), .QN(n337) );
  AO22X1 U462 ( .IN1(n322), .IN2(n321), .IN3(n319), .IN4(n58), .Q(n338) );
  XOR2X1 U463 ( .IN1(g471), .IN2(n806), .Q(n319) );
  XOR2X1 U464 ( .IN1(n340), .IN2(g471), .Q(n321) );
  NAND4X0 U465 ( .IN1(g206), .IN2(n343), .IN3(n344), .IN4(n345), .QN(n342) );
  OR2X1 U467 ( .IN1(n346), .IN2(g690), .Q(n344) );
  NAND3X0 U469 ( .IN1(n347), .IN2(n75), .IN3(n348), .QN(n341) );
  OA22X1 U470 ( .IN1(n787), .IN2(n349), .IN3(g694), .IN4(n346), .Q(n348) );
  NAND4X0 U473 ( .IN1(n352), .IN2(n866), .IN3(n351), .IN4(n350), .QN(g6485) );
  AOI221X1 U474 ( .IN1(g5629), .IN2(n876), .IN3(g5630), .IN4(n979), .IN5(n353), 
        .QN(n352) );
  NAND4X0 U477 ( .IN1(n354), .IN2(n866), .IN3(n355), .IN4(n356), .QN(g6483) );
  AOI221X1 U478 ( .IN1(g5533), .IN2(n974), .IN3(n979), .IN4(g5535), .IN5(n357), 
        .QN(n356) );
  AOI221X1 U482 ( .IN1(g561), .IN2(n962), .IN3(n953), .IN4(n1035), .IN5(n3), 
        .QN(n361) );
  AOI221X1 U487 ( .IN1(g562), .IN2(n962), .IN3(n756), .IN4(n955), .IN5(n3), 
        .QN(n368) );
  AOI221X1 U492 ( .IN1(g672), .IN2(n374), .IN3(g563), .IN4(n962), .IN5(n375), 
        .QN(n373) );
  OA221X1 U495 ( .IN1(n376), .IN2(n108), .IN3(n770), .IN4(n96), .IN5(n377), 
        .Q(n371) );
  OA22X1 U496 ( .IN1(g489), .IN2(n378), .IN3(n379), .IN4(n81), .Q(n377) );
  AOI221X1 U499 ( .IN1(g669), .IN2(n374), .IN3(g564), .IN4(n961), .IN5(n384), 
        .QN(n383) );
  AND4X1 U501 ( .IN1(n387), .IN2(n770), .IN3(n378), .IN4(n376), .Q(n386) );
  AND4X1 U509 ( .IN1(n4), .IN2(n104), .IN3(g680), .IN4(n393), .Q(n374) );
  OA221X1 U514 ( .IN1(n376), .IN2(n44), .IN3(n770), .IN4(n122), .IN5(n399), 
        .Q(n381) );
  OA22X1 U515 ( .IN1(g486), .IN2(n378), .IN3(n956), .IN4(n18), .Q(n399) );
  NOR3X0 U520 ( .IN1(n991), .IN2(g680), .IN3(n395), .QN(n392) );
  NAND4X0 U525 ( .IN1(n400), .IN2(g699), .IN3(n1027), .IN4(g702), .QN(n394) );
  AO21X1 U526 ( .IN1(g266), .IN2(n1038), .IN3(n265), .Q(n400) );
  AND2X1 U531 ( .IN1(g662), .IN2(n1038), .Q(n265) );
  AO21X1 U535 ( .IN1(n767), .IN2(n410), .IN3(n741), .Q(g6455) );
  AO21X1 U539 ( .IN1(n417), .IN2(n786), .IN3(n1023), .Q(g6454) );
  AO21X1 U542 ( .IN1(n767), .IN2(n424), .IN3(n1025), .Q(g6453) );
  XOR2X1 U543 ( .IN1(g69), .IN2(n425), .Q(n424) );
  AO21X1 U546 ( .IN1(n429), .IN2(n786), .IN3(n1023), .Q(g6452) );
  AO21X1 U549 ( .IN1(n767), .IN2(n432), .IN3(n1025), .Q(g6450) );
  XOR2X1 U550 ( .IN1(n137), .IN2(n433), .Q(n432) );
  OR2X1 U552 ( .IN1(n437), .IN2(g54), .Q(n420) );
  AO21X1 U553 ( .IN1(n786), .IN2(n438), .IN3(n741), .Q(g6447) );
  NAND4X0 U556 ( .IN1(g49), .IN2(g361), .IN3(n1013), .IN4(n719), .QN(n436) );
  NAND4X0 U557 ( .IN1(n774), .IN2(n1013), .IN3(n55), .IN4(n132), .QN(n437) );
  OAI21X1 U560 ( .IN1(n446), .IN2(n894), .IN3(g49), .QN(n444) );
  AO22X1 U561 ( .IN1(g370), .IN2(n407), .IN3(n448), .IN4(n707), .Q(n447) );
  XOR2X1 U562 ( .IN1(g361), .IN2(n774), .Q(n448) );
  NAND3X0 U567 ( .IN1(n455), .IN2(n154), .IN3(n147), .QN(n241) );
  AOI22X1 U569 ( .IN1(n408), .IN2(g84), .IN3(n409), .IN4(n28), .QN(n460) );
  NAND4X0 U571 ( .IN1(n423), .IN2(n55), .IN3(n461), .IN4(n132), .QN(n416) );
  OAI21X1 U576 ( .IN1(n8), .IN2(n1014), .IN3(n456), .QN(n464) );
  AO22X1 U588 ( .IN1(n21), .IN2(n953), .IN3(g297), .IN4(n708), .Q(g6298) );
  AO22X1 U592 ( .IN1(n21), .IN2(n955), .IN3(g293), .IN4(n708), .Q(g6294) );
  AO22X1 U593 ( .IN1(n20), .IN2(n955), .IN3(n478), .IN4(g536), .Q(g6293) );
  AO22X1 U595 ( .IN1(n881), .IN2(n981), .IN3(g500), .IN4(n975), .Q(g6292) );
  AO21X1 U597 ( .IN1(n466), .IN2(g594), .IN3(n159), .Q(n474) );
  AND2X1 U598 ( .IN1(g582), .IN2(n477), .Q(n473) );
  AND2X1 U599 ( .IN1(n877), .IN2(n848), .Q(n477) );
  AND2X1 U609 ( .IN1(n489), .IN2(n490), .Q(g6142) );
  NAND4X0 U610 ( .IN1(n115), .IN2(g594), .IN3(n491), .IN4(g574), .QN(n490) );
  NAND3X0 U611 ( .IN1(n492), .IN2(n493), .IN3(n494), .QN(n489) );
  XOR2X1 U612 ( .IN1(n777), .IN2(g594), .Q(n494) );
  NAND4X0 U613 ( .IN1(g586), .IN2(n495), .IN3(n496), .IN4(n497), .QN(n493) );
  NAND3X0 U616 ( .IN1(n499), .IN2(n89), .IN3(n500), .QN(n492) );
  OA22X1 U617 ( .IN1(g582), .IN2(n501), .IN3(n842), .IN4(n498), .Q(n500) );
  OA22X1 U618 ( .IN1(n898), .IN2(g578), .IN3(n846), .IN4(n116), .Q(n501) );
  AO21X1 U620 ( .IN1(n502), .IN2(n503), .IN3(n890), .Q(g6118) );
  XOR2X1 U621 ( .IN1(g188), .IN2(n504), .Q(n503) );
  OA221X1 U622 ( .IN1(g193), .IN2(n950), .IN3(n505), .IN4(n506), .IN5(n969), 
        .Q(n504) );
  OA221X1 U625 ( .IN1(g184), .IN2(n951), .IN3(n505), .IN4(n512), .IN5(n970), 
        .Q(n511) );
  AO21X1 U631 ( .IN1(n502), .IN2(n518), .IN3(n682), .Q(g6113) );
  XOR2X1 U632 ( .IN1(g161), .IN2(n520), .Q(n518) );
  OA221X1 U633 ( .IN1(g166), .IN2(n950), .IN3(n505), .IN4(n521), .IN5(n969), 
        .Q(n520) );
  XOR3X1 U634 ( .IN1(n524), .IN2(n525), .IN3(n526), .Q(g6658) );
  XOR3X1 U635 ( .IN1(g6686), .IN2(g6685), .IN3(n527), .Q(n526) );
  XOR2X1 U636 ( .IN1(n84), .IN2(g6688), .Q(n527) );
  XOR2X1 U637 ( .IN1(g6690), .IN2(g6689), .Q(n525) );
  XOR2X1 U638 ( .IN1(g6684), .IN2(g6691), .Q(n524) );
  AO21X1 U641 ( .IN1(n38), .IN2(n969), .IN3(n133), .Q(n529) );
  AO22X1 U642 ( .IN1(g157), .IN2(n505), .IN3(n533), .IN4(n950), .Q(n532) );
  AO21X1 U646 ( .IN1(n37), .IN2(n970), .IN3(n106), .Q(n536) );
  OR2X1 U647 ( .IN1(n951), .IN2(g148), .Q(n539) );
  AO221X1 U650 ( .IN1(g366), .IN2(n545), .IN3(g398), .IN4(n987), .IN5(n749), 
        .Q(g5916) );
  OA221X1 U651 ( .IN1(n546), .IN2(g111), .IN3(n125), .IN4(n547), .IN5(n827), 
        .Q(g5701) );
  OA22X1 U653 ( .IN1(n51), .IN2(n509), .IN3(g188), .IN4(n508), .Q(n548) );
  NAND3X0 U654 ( .IN1(n513), .IN2(n45), .IN3(n109), .QN(n508) );
  OAI21X1 U659 ( .IN1(n11), .IN2(n541), .IN3(n543), .QN(n549) );
  AO22X1 U661 ( .IN1(g394), .IN2(n69), .IN3(n915), .IN4(g398), .Q(g5700) );
  AO22X1 U662 ( .IN1(n987), .IN2(g390), .IN3(g394), .IN4(n914), .Q(g5699) );
  AO22X1 U663 ( .IN1(n987), .IN2(g386), .IN3(n915), .IN4(g390), .Q(g5698) );
  AO22X1 U664 ( .IN1(n987), .IN2(g382), .IN3(n916), .IN4(g386), .Q(g5697) );
  AO22X1 U665 ( .IN1(n987), .IN2(g378), .IN3(n915), .IN4(g382), .Q(g5696) );
  AO22X1 U666 ( .IN1(n69), .IN2(g374), .IN3(n916), .IN4(g378), .Q(g5695) );
  AO22X1 U667 ( .IN1(n987), .IN2(g370), .IN3(n914), .IN4(g374), .Q(g5694) );
  AO22X1 U668 ( .IN1(n69), .IN2(g366), .IN3(n916), .IN4(g370), .Q(g5693) );
  AO22X1 U670 ( .IN1(n739), .IN2(n1011), .IN3(n551), .IN4(n32), .Q(g5630) );
  AO22X1 U672 ( .IN1(n739), .IN2(n1016), .IN3(n554), .IN4(n13), .Q(g5629) );
  AO22X1 U675 ( .IN1(n955), .IN2(n1039), .IN3(n563), .IN4(n562), .Q(g5627) );
  AOI21X1 U676 ( .IN1(n917), .IN2(n34), .IN3(n560), .QN(n562) );
  AO22X1 U678 ( .IN1(n875), .IN2(n1011), .IN3(n563), .IN4(n569), .Q(g5625) );
  AOI21X1 U680 ( .IN1(n346), .IN2(n75), .IN3(n789), .QN(n570) );
  AO22X1 U681 ( .IN1(g691), .IN2(n1009), .IN3(n572), .IN4(n571), .Q(g5622) );
  AO221X1 U682 ( .IN1(g148), .IN2(n573), .IN3(g193), .IN4(n807), .IN5(n140), 
        .Q(g5583) );
  NAND3X0 U684 ( .IN1(n575), .IN2(n31), .IN3(n32), .QN(n574) );
  NAND3X0 U687 ( .IN1(n577), .IN2(n12), .IN3(n13), .QN(n576) );
  XOR2X1 U693 ( .IN1(n113), .IN2(g281), .Q(n311) );
  NOR3X0 U694 ( .IN1(g283), .IN2(g478), .IN3(g282), .QN(n578) );
  AO21X1 U697 ( .IN1(n806), .IN2(n579), .IN3(n14), .Q(n566) );
  XOR2X1 U699 ( .IN1(n59), .IN2(g209), .Q(n322) );
  NOR3X0 U700 ( .IN1(g211), .IN2(g471), .IN3(g210), .QN(n579) );
  AO22X1 U701 ( .IN1(g184), .IN2(n807), .IN3(n580), .IN4(g193), .Q(g5474) );
  AO22X1 U702 ( .IN1(g175), .IN2(n807), .IN3(g184), .IN4(n580), .Q(g5473) );
  AO22X1 U703 ( .IN1(g166), .IN2(n807), .IN3(g175), .IN4(n580), .Q(g5472) );
  AO22X1 U704 ( .IN1(n807), .IN2(g157), .IN3(g166), .IN4(n580), .Q(g5471) );
  AO22X1 U705 ( .IN1(n807), .IN2(g148), .IN3(n580), .IN4(g157), .Q(g5470) );
  AO21X1 U707 ( .IN1(n162), .IN2(n144), .IN3(g669), .Q(g5386) );
  XOR2X1 U710 ( .IN1(g4101), .IN2(g4100), .Q(n584) );
  XOR2X1 U711 ( .IN1(g4103), .IN2(g4102), .Q(n582) );
  AO21X1 U715 ( .IN1(g357), .IN2(n588), .IN3(n68), .Q(g5303) );
  AO221X1 U717 ( .IN1(n590), .IN2(n66), .IN3(g349), .IN4(n591), .IN5(n68), .Q(
        g5295) );
  AO221X1 U719 ( .IN1(n704), .IN2(n594), .IN3(n66), .IN4(n595), .IN5(n68), .Q(
        g5291) );
  OR2X1 U720 ( .IN1(n595), .IN2(n71), .Q(n594) );
  NAND3X0 U721 ( .IN1(n597), .IN2(n596), .IN3(n826), .QN(g5277) );
  OAI21X1 U722 ( .IN1(n71), .IN2(n706), .IN3(g341), .QN(n597) );
  AND2X1 U734 ( .IN1(n589), .IN2(g323), .Q(n609) );
  NOR3X0 U736 ( .IN1(n111), .IN2(n606), .IN3(n610), .QN(g5017) );
  AND2X1 U737 ( .IN1(n611), .IN2(g654), .Q(n606) );
  AND2X1 U739 ( .IN1(g628), .IN2(n613), .Q(n604) );
  XOR2X1 U740 ( .IN1(g128), .IN2(n124), .Q(n614) );
  NOR3X0 U741 ( .IN1(n111), .IN2(n611), .IN3(n615), .QN(g4761) );
  AND2X1 U742 ( .IN1(n616), .IN2(g650), .Q(n611) );
  AO21X1 U743 ( .IN1(g139), .IN2(n617), .IN3(n35), .Q(g4757) );
  AO221X1 U745 ( .IN1(g135), .IN2(n619), .IN3(n40), .IN4(n620), .IN5(n35), .Q(
        g4752) );
  OR2X1 U746 ( .IN1(n620), .IN2(n124), .Q(n619) );
  OAI21X1 U750 ( .IN1(n124), .IN2(g128), .IN3(g131), .QN(n622) );
  NOR3X0 U753 ( .IN1(n111), .IN2(n616), .IN3(n626), .QN(g4501) );
  AND2X1 U754 ( .IN1(n627), .IN2(g646), .Q(n616) );
  AND2X1 U756 ( .IN1(n630), .IN2(g622), .Q(n624) );
  AO22X1 U757 ( .IN1(n802), .IN2(g422), .IN3(g426), .IN4(n1034), .Q(g4458) );
  AO22X1 U758 ( .IN1(n1043), .IN2(g418), .IN3(g422), .IN4(n1033), .Q(g4455) );
  AO22X1 U759 ( .IN1(n802), .IN2(g449), .IN3(g445), .IN4(n1034), .Q(g4454) );
  AO22X1 U760 ( .IN1(n1042), .IN2(g414), .IN3(g418), .IN4(n1033), .Q(g4451) );
  AO22X1 U761 ( .IN1(n1043), .IN2(g453), .IN3(g449), .IN4(n1034), .Q(g4450) );
  AO22X1 U762 ( .IN1(n1042), .IN2(g410), .IN3(g414), .IN4(n1033), .Q(g4447) );
  AO22X1 U763 ( .IN1(n802), .IN2(g457), .IN3(g453), .IN4(n1034), .Q(g4446) );
  AO22X1 U764 ( .IN1(n1042), .IN2(g406), .IN3(g410), .IN4(n1033), .Q(g4444) );
  AO22X1 U765 ( .IN1(n1043), .IN2(g461), .IN3(g457), .IN4(n1034), .Q(g4443) );
  AO22X1 U766 ( .IN1(n1042), .IN2(g402), .IN3(g406), .IN4(n1033), .Q(g4441) );
  AO22X1 U767 ( .IN1(n802), .IN2(g430), .IN3(g461), .IN4(n1034), .Q(g4440) );
  AO22X1 U769 ( .IN1(g465), .IN2(g478), .IN3(g471), .IN4(n27), .Q(n632) );
  AO22X1 U770 ( .IN1(n1042), .IN2(g437), .IN3(g434), .IN4(n1032), .Q(g4436) );
  AO22X1 U771 ( .IN1(n1043), .IN2(g426), .IN3(g430), .IN4(n1032), .Q(g4434) );
  AO22X1 U772 ( .IN1(n1042), .IN2(g441), .IN3(g437), .IN4(n1032), .Q(g4433) );
  AO22X1 U773 ( .IN1(n802), .IN2(g445), .IN3(g441), .IN4(n1032), .Q(g4430) );
  XOR2X1 U777 ( .IN1(g528), .IN2(g254), .Q(n639) );
  XOR2X1 U778 ( .IN1(g524), .IN2(g248), .Q(n638) );
  XOR2X1 U779 ( .IN1(g520), .IN2(g242), .Q(n637) );
  NOR3X0 U780 ( .IN1(n641), .IN2(n642), .IN3(n643), .QN(n635) );
  XOR2X1 U781 ( .IN1(g500), .IN2(g212), .Q(n643) );
  XOR2X1 U782 ( .IN1(g508), .IN2(g224), .Q(n642) );
  XOR2X1 U783 ( .IN1(g504), .IN2(g218), .Q(n641) );
  XNOR2X1 U784 ( .IN1(g230), .IN2(g512), .Q(n634) );
  XNOR2X1 U785 ( .IN1(g236), .IN2(g516), .Q(n633) );
  NOR3X0 U786 ( .IN1(n766), .IN2(n627), .IN3(n644), .QN(g4219) );
  AND2X1 U787 ( .IN1(n645), .IN2(g606), .Q(n627) );
  NOR3X0 U790 ( .IN1(n766), .IN2(n645), .IN3(n648), .QN(g3844) );
  AND2X1 U795 ( .IN1(g331), .IN2(n625), .Q(g3731) );
  AND2X1 U796 ( .IN1(n625), .IN2(g328), .Q(g3730) );
  AND2X1 U797 ( .IN1(g327), .IN2(n625), .Q(g3729) );
  AND2X1 U798 ( .IN1(g326), .IN2(n625), .Q(g3728) );
  AND2X1 U801 ( .IN1(g122), .IN2(n628), .Q(g3727) );
  AND2X1 U802 ( .IN1(n628), .IN2(g119), .Q(g3726) );
  AND2X1 U803 ( .IN1(g118), .IN2(n628), .Q(g3725) );
  AND2X1 U804 ( .IN1(g117), .IN2(n628), .Q(g3724) );
  AND2X1 U806 ( .IN1(n189), .IN2(n193), .Q(n542) );
  OA22X1 U809 ( .IN1(g3599), .IN2(n42), .IN3(n76), .IN4(n111), .Q(n653) );
  AND2X1 U810 ( .IN1(g634), .IN2(n219), .Q(n214) );
  NOR3X0 U811 ( .IN1(n766), .IN2(n219), .IN3(n213), .QN(g2859) );
  OA22X1 U814 ( .IN1(g489), .IN2(n108), .IN3(g486), .IN4(n44), .Q(g2433) );
  INVX0 U816 ( .INP(1'b1), .ZN(g6728) );
  INVX0 U818 ( .INP(1'b1), .ZN(g5692) );
  NOR2X1 U820 ( .IN1(n693), .IN2(n692), .QN(n408) );
  DELLN2X2 U821 ( .INP(g14), .Z(n815) );
  IBUFFX16 U822 ( .INP(n397), .ZN(n911) );
  AND3X1 U823 ( .IN1(n397), .IN2(g683), .IN3(n86), .Q(n886) );
  INVX1 U824 ( .INP(n891), .ZN(n892) );
  NOR4X1 U825 ( .IN1(n973), .IN2(n847), .IN3(n972), .IN4(n957), .QN(n387) );
  DELLN1X2 U826 ( .INP(n401), .Z(n737) );
  AO21X1 U827 ( .IN1(n844), .IN2(n578), .IN3(n33), .Q(n559) );
  NOR3X0 U828 ( .IN1(g689), .IN2(g698), .IN3(g688), .QN(n263) );
  INVX0 U829 ( .INP(n788), .ZN(n458) );
  AND3X1 U830 ( .IN1(n840), .IN2(n397), .IN3(n264), .Q(n487) );
  NAND3X0 U831 ( .IN1(n396), .IN2(g677), .IN3(n398), .QN(n369) );
  NBUFFX2 U832 ( .INP(n309), .Z(n860) );
  NAND3X0 U833 ( .IN1(n4), .IN2(n104), .IN3(n851), .QN(n376) );
  NAND3X0 U834 ( .IN1(n396), .IN2(n128), .IN3(n398), .QN(n362) );
  NAND3X0 U835 ( .IN1(n264), .IN2(n100), .IN3(n912), .QN(n475) );
  NAND3X1 U836 ( .IN1(g64), .IN2(g59), .IN3(g69), .QN(n421) );
  AND2X1 U837 ( .IN1(g625), .IN2(n624), .Q(n613) );
  INVX0 U838 ( .INP(n416), .ZN(n54) );
  AND2X1 U839 ( .IN1(n877), .IN2(n878), .Q(n674) );
  NBUFFX2 U840 ( .INP(n14), .Z(n852) );
  NBUFFX2 U841 ( .INP(n973), .Z(n876) );
  NAND3X0 U842 ( .IN1(n843), .IN2(n203), .IN3(n171), .QN(n195) );
  OAI21X1 U843 ( .IN1(n864), .IN2(n859), .IN3(n753), .QN(g6456) );
  NOR3X0 U844 ( .IN1(n870), .IN2(n624), .IN3(n629), .QN(g4460) );
  DELLN1X2 U845 ( .INP(g18), .Z(n812) );
  NBUFFX2 U846 ( .INP(g24), .Z(n818) );
  AO22X1 U847 ( .IN1(g545), .IN2(n959), .IN3(n960), .IN4(n230), .Q(g6787) );
  DELLN1X2 U848 ( .INP(g10), .Z(n816) );
  NBUFFX2 U849 ( .INP(n771), .Z(n801) );
  AO22X1 U850 ( .IN1(n1039), .IN2(n842), .IN3(n992), .IN4(n574), .Q(g5535) );
  OR2X1 U851 ( .IN1(g610), .IN2(g602), .Q(n654) );
  DELLN1X2 U852 ( .INP(g1), .Z(n817) );
  DELLN1X2 U853 ( .INP(g6), .Z(n823) );
  DELLN1X2 U854 ( .INP(g2), .Z(n824) );
  AND2X1 U855 ( .IN1(n263), .IN2(n94), .Q(n662) );
  NBUFFX2 U856 ( .INP(n415), .Z(n719) );
  NAND2X1 U857 ( .IN1(n462), .IN2(n459), .QN(n415) );
  AO21X1 U858 ( .IN1(n113), .IN2(n561), .IN3(n553), .Q(n575) );
  DELLN1X2 U859 ( .INP(n553), .Z(n677) );
  AND2X1 U860 ( .IN1(g278), .IN2(n828), .Q(n560) );
  NAND2X0 U861 ( .IN1(g207), .IN2(n567), .QN(n568) );
  AO22X2 U862 ( .IN1(n1036), .IN2(g682), .IN3(n989), .IN4(n280), .Q(n275) );
  DELLN1X2 U863 ( .INP(n409), .Z(n699) );
  NAND2X1 U864 ( .IN1(n385), .IN2(n386), .QN(n284) );
  NAND3X0 U865 ( .IN1(n389), .IN2(n750), .IN3(n843), .QN(n756) );
  NAND3X0 U866 ( .IN1(n202), .IN2(n172), .IN3(n389), .QN(n291) );
  NAND2X1 U867 ( .IN1(n664), .IN2(n784), .QN(n663) );
  AO22X2 U868 ( .IN1(n898), .IN2(n1009), .IN3(n990), .IN4(n759), .Q(g6792) );
  AO221X2 U869 ( .IN1(n275), .IN2(g683), .IN3(n276), .IN4(g685), .IN5(n990), 
        .Q(n274) );
  NAND2X1 U870 ( .IN1(n712), .IN2(n662), .QN(n838) );
  INVX0 U871 ( .INP(n838), .ZN(n974) );
  NBUFFX2 U872 ( .INP(n586), .Z(n771) );
  DELLN1X2 U873 ( .INP(n86), .Z(n1029) );
  XOR2X2 U874 ( .IN1(n72), .IN2(g291), .Q(n227) );
  NOR3X2 U875 ( .IN1(g685), .IN2(g688), .IN3(n391), .QN(n174) );
  NOR2X0 U876 ( .IN1(n663), .IN2(n291), .QN(n385) );
  NOR2X0 U877 ( .IN1(n961), .IN2(n374), .QN(n664) );
  NBUFFX2 U878 ( .INP(n291), .Z(n1035) );
  NAND3X1 U879 ( .IN1(n165), .IN2(n160), .IN3(g107), .QN(n573) );
  NOR4X0 U880 ( .IN1(n72), .IN2(n57), .IN3(n391), .IN4(g688), .QN(n397) );
  INVX0 U881 ( .INP(n982), .ZN(n880) );
  NAND3X0 U882 ( .IN1(n392), .IN2(g679), .IN3(g678), .QN(n927) );
  NOR2X0 U883 ( .IN1(n906), .IN2(n908), .QN(n567) );
  NBUFFX2 U884 ( .INP(n1015), .Z(n721) );
  OR2X1 U885 ( .IN1(n105), .IN2(n925), .Q(n924) );
  NBUFFX2 U886 ( .INP(n1037), .Z(n1031) );
  NAND3X0 U887 ( .IN1(n886), .IN2(n48), .IN3(g681), .QN(n364) );
  AND3X1 U888 ( .IN1(n456), .IN2(n457), .IN3(n235), .Q(n780) );
  AND2X1 U889 ( .IN1(n783), .IN2(n827), .Q(n747) );
  NBUFFX2 U890 ( .INP(n721), .Z(n1026) );
  DELLN1X2 U891 ( .INP(n630), .Z(n893) );
  NBUFFX2 U892 ( .INP(n567), .Z(n789) );
  INVX0 U893 ( .INP(n468), .ZN(n778) );
  INVX0 U894 ( .INP(n723), .ZN(n593) );
  INVX0 U895 ( .INP(n751), .ZN(n752) );
  INVX0 U896 ( .INP(n713), .ZN(n407) );
  INVX0 U897 ( .INP(n959), .ZN(n960) );
  NBUFFX2 U898 ( .INP(n473), .Z(n799) );
  NBUFFX2 U899 ( .INP(n182), .Z(n827) );
  INVX0 U900 ( .INP(n182), .ZN(n140) );
  NAND3X0 U901 ( .IN1(n174), .IN2(n793), .IN3(n175), .QN(n203) );
  XNOR2X1 U902 ( .IN1(n898), .IN2(n191), .Q(n184) );
  NBUFFX2 U903 ( .INP(n522), .Z(n820) );
  NBUFFX2 U904 ( .INP(n471), .Z(n748) );
  AO22X1 U905 ( .IN1(n20), .IN2(n875), .IN3(g465), .IN4(n748), .Q(g6297) );
  AOI222X1 U906 ( .IN1(g5531), .IN2(n974), .IN3(n865), .IN4(g402), .IN5(g5532), 
        .IN6(n679), .QN(n380) );
  NOR3X0 U907 ( .IN1(n677), .IN2(g281), .IN3(n918), .QN(n552) );
  AO22X1 U908 ( .IN1(n881), .IN2(n842), .IN3(g516), .IN4(n716), .Q(g6307) );
  NOR3X0 U909 ( .IN1(n809), .IN2(g209), .IN3(n909), .QN(n555) );
  XOR2X1 U910 ( .IN1(g532), .IN2(g260), .Q(n640) );
  AOI22X1 U911 ( .IN1(g571), .IN2(n1031), .IN3(g260), .IN4(n983), .QN(n266) );
  AO22X1 U912 ( .IN1(n986), .IN2(n968), .IN3(g212), .IN4(n880), .Q(n255) );
  NAND3X1 U913 ( .IN1(n396), .IN2(g682), .IN3(g677), .QN(n715) );
  NBUFFX2 U914 ( .INP(n87), .Z(n1041) );
  XOR2X1 U915 ( .IN1(g684), .IN2(g290), .Q(n228) );
  AND2X1 U916 ( .IN1(g606), .IN2(n198), .Q(n201) );
  AO22X1 U917 ( .IN1(g678), .IN2(n983), .IN3(g642), .IN4(n967), .Q(n198) );
  AND2X1 U918 ( .IN1(n398), .IN2(g683), .Q(n840) );
  OA22X1 U919 ( .IN1(g697), .IN2(n754), .IN3(g696), .IN4(n119), .Q(n349) );
  NAND3X1 U920 ( .IN1(n119), .IN2(n17), .IN3(g205), .QN(n347) );
  AO221X1 U921 ( .IN1(g693), .IN2(n760), .IN3(g692), .IN4(n754), .IN5(n787), 
        .Q(n343) );
  NBUFFX2 U922 ( .INP(n913), .Z(n790) );
  NBUFFX2 U923 ( .INP(n1041), .Z(n993) );
  OAI22X1 U924 ( .IN1(n266), .IN2(n993), .IN3(n772), .IN4(n110), .QN(n1006) );
  AO22X1 U925 ( .IN1(n965), .IN2(n1031), .IN3(g218), .IN4(n880), .Q(n250) );
  AO22X1 U926 ( .IN1(g680), .IN2(n1039), .IN3(g269), .IN4(n256), .Q(n251) );
  AO22X1 U927 ( .IN1(g678), .IN2(n993), .IN3(g269), .IN4(n255), .Q(n249) );
  AO22X1 U928 ( .IN1(g654), .IN2(n968), .IN3(g254), .IN4(n880), .Q(n278) );
  NBUFFX2 U929 ( .INP(n87), .Z(n1039) );
  AND3X1 U930 ( .IN1(n192), .IN2(n190), .IN3(n680), .Q(n167) );
  NAND3X0 U931 ( .IN1(g678), .IN2(n104), .IN3(n851), .QN(n378) );
  INVX0 U932 ( .INP(n698), .ZN(n188) );
  DELLN1X2 U933 ( .INP(n781), .Z(n698) );
  AND2X1 U934 ( .IN1(n160), .IN2(n192), .Q(n187) );
  NAND3X0 U935 ( .IN1(n171), .IN2(n173), .IN3(n750), .QN(n169) );
  NAND3X0 U936 ( .IN1(n755), .IN2(n174), .IN3(n175), .QN(n173) );
  DELLN1X2 U937 ( .INP(n568), .Z(n849) );
  INVX0 U938 ( .INP(g532), .ZN(n135) );
  NAND3X0 U939 ( .IN1(n116), .IN2(n136), .IN3(g582), .QN(n497) );
  NAND3X0 U940 ( .IN1(n116), .IN2(n17), .IN3(g582), .QN(n499) );
  XNOR3X1 U941 ( .IN1(n584), .IN2(g4099), .IN3(n744), .Q(n933) );
  OR2X1 U942 ( .IN1(n695), .IN2(g64), .Q(n427) );
  AOI22X1 U943 ( .IN1(g557), .IN2(n961), .IN3(g528), .IN4(n24), .QN(n285) );
  INVX0 U944 ( .INP(n763), .ZN(n802) );
  INVX0 U945 ( .INP(n423), .ZN(n80) );
  NBUFFX2 U946 ( .INP(n707), .Z(n1012) );
  INVX0 U947 ( .INP(g209), .ZN(n114) );
  AO22X1 U948 ( .IN1(g682), .IN2(n993), .IN3(n772), .IN4(n280), .Q(n281) );
  INVX0 U949 ( .INP(g613), .ZN(n105) );
  AND2X1 U950 ( .IN1(g642), .IN2(g634), .Q(n814) );
  INVX0 U951 ( .INP(n556), .ZN(n808) );
  NBUFFX2 U952 ( .INP(n700), .Z(n922) );
  INVX0 U953 ( .INP(n837), .ZN(n301) );
  NAND3X0 U954 ( .IN1(n888), .IN2(n143), .IN3(n697), .QN(n543) );
  AO222X1 U955 ( .IN1(g5622), .IN2(n974), .IN3(n865), .IN4(g406), .IN5(g5625), 
        .IN6(n978), .Q(n718) );
  INVX0 U956 ( .INP(n631), .ZN(n1042) );
  XOR2X1 U957 ( .IN1(n795), .IN2(g143), .Q(n533) );
  NBUFFX2 U958 ( .INP(n333), .Z(n917) );
  INVX0 U959 ( .INP(n845), .ZN(n502) );
  INVX0 U960 ( .INP(n930), .ZN(n975) );
  INVX0 U961 ( .INP(n155), .ZN(g4110) );
  OR2X1 U962 ( .IN1(g337), .IN2(n171), .Q(n296) );
  OAI21X1 U963 ( .IN1(n884), .IN2(n871), .IN3(n519), .QN(g6116) );
  NAND3X0 U964 ( .IN1(n685), .IN2(n452), .IN3(n453), .QN(n451) );
  NOR3X0 U965 ( .IN1(n159), .IN2(n893), .IN3(n646), .QN(g4157) );
  AO22X1 U966 ( .IN1(n955), .IN2(n1009), .IN3(n570), .IN4(n571), .Q(g5624) );
  AO22X1 U967 ( .IN1(n881), .IN2(n898), .IN3(g528), .IN4(n975), .Q(g6286) );
  AO22X1 U968 ( .IN1(g402), .IN2(n1033), .IN3(n1043), .IN4(n632), .Q(g4438) );
  AO22X1 U969 ( .IN1(n21), .IN2(n875), .IN3(n992), .IN4(n475), .Q(g6290) );
  AND3X1 U970 ( .IN1(n593), .IN2(n103), .IN3(g349), .Q(n592) );
  AND2X1 U971 ( .IN1(n472), .IN2(n779), .Q(n800) );
  NOR2X0 U972 ( .IN1(n605), .IN2(n766), .QN(g5149) );
  XNOR2X1 U973 ( .IN1(n606), .IN2(g571), .Q(n605) );
  AOI22X1 U974 ( .IN1(g558), .IN2(n962), .IN3(g524), .IN4(n861), .QN(n293) );
  NAND3X1 U975 ( .IN1(n589), .IN2(n101), .IN3(g323), .QN(n588) );
  AO22X1 U976 ( .IN1(n882), .IN2(n875), .IN3(g504), .IN4(n975), .Q(g6296) );
  AO22X1 U977 ( .IN1(n20), .IN2(n953), .IN3(n484), .IN4(n748), .Q(g6289) );
  AO22X1 U978 ( .IN1(n852), .IN2(n27), .IN3(g465), .IN4(n857), .Q(n486) );
  XOR2X1 U979 ( .IN1(n706), .IN2(n71), .Q(n587) );
  INVX0 U980 ( .INP(n722), .ZN(n67) );
  OR2X1 U981 ( .IN1(n682), .IN2(n858), .Q(g6108) );
  NAND3X0 U982 ( .IN1(n538), .IN2(n970), .IN3(n539), .QN(n537) );
  AND2X1 U983 ( .IN1(n919), .IN2(n441), .Q(n929) );
  OA22X1 U984 ( .IN1(n774), .IN2(n414), .IN3(n54), .IN4(n719), .Q(n412) );
  NAND3X0 U985 ( .IN1(n618), .IN2(n129), .IN3(g114), .QN(n617) );
  AOI22X1 U986 ( .IN1(g559), .IN2(n962), .IN3(g520), .IN4(n861), .QN(n351) );
  AO22X1 U987 ( .IN1(n981), .IN2(n1017), .IN3(n571), .IN4(n760), .Q(g5531) );
  AO22X1 U988 ( .IN1(n882), .IN2(n955), .IN3(g508), .IN4(n716), .Q(g6300) );
  AO22X1 U989 ( .IN1(n882), .IN2(n846), .IN3(g524), .IN4(n975), .Q(g6310) );
  NAND3X0 U990 ( .IN1(n622), .IN2(n834), .IN3(n166), .QN(g4740) );
  AOI22X1 U991 ( .IN1(g560), .IN2(n962), .IN3(g516), .IN4(n861), .QN(n355) );
  NAND3X0 U992 ( .IN1(n446), .IN2(n447), .IN3(n685), .QN(n445) );
  INVX0 U993 ( .INP(n193), .ZN(n139) );
  AO22X1 U994 ( .IN1(n882), .IN2(n953), .IN3(g512), .IN4(n975), .Q(g6303) );
  AO22X1 U995 ( .IN1(n20), .IN2(n981), .IN3(g532), .IN4(n748), .Q(g6301) );
  INVX0 U996 ( .INP(n879), .ZN(n968) );
  NAND3X0 U997 ( .IN1(n721), .IN2(n703), .IN3(g319), .QN(n545) );
  OR2X1 U998 ( .IN1(g64), .IN2(g69), .Q(n665) );
  AND2X1 U999 ( .IN1(n195), .IN2(n170), .Q(n666) );
  AND2X1 U1000 ( .IN1(n540), .IN2(n773), .Q(n839) );
  OR2X1 U1001 ( .IN1(n416), .IN2(g79), .Q(n667) );
  AND2X1 U1002 ( .IN1(n382), .IN2(n381), .Q(n668) );
  OR2X1 U1003 ( .IN1(n114), .IN2(g208), .Q(n669) );
  AND3X1 U1004 ( .IN1(n238), .IN2(g328), .IN3(n239), .Q(n670) );
  AND2X1 U1005 ( .IN1(n106), .IN2(n133), .Q(n671) );
  AND2X1 U1006 ( .IN1(n901), .IN2(n900), .Q(n672) );
  AND3X1 U1007 ( .IN1(n285), .IN2(n283), .IN3(n910), .Q(n673) );
  AND2X1 U1008 ( .IN1(g179), .IN2(g170), .Q(n675) );
  AND3X1 U1009 ( .IN1(g152), .IN2(n675), .IN3(g143), .Q(n676) );
  INVX0 U1010 ( .INP(n982), .ZN(n983) );
  INVX0 U1011 ( .INP(g84), .ZN(n28) );
  NOR3X0 U1012 ( .IN1(n740), .IN2(n477), .IN3(n482), .QN(g6291) );
  NBUFFX2 U1013 ( .INP(n304), .Z(n678) );
  NBUFFX2 U1014 ( .INP(n978), .Z(n679) );
  NBUFFX2 U1015 ( .INP(n542), .Z(n680) );
  NAND3X0 U1016 ( .IN1(n152), .IN2(n913), .IN3(n684), .QN(n459) );
  OR2X1 U1017 ( .IN1(n161), .IN2(n757), .Q(n189) );
  INVX0 U1018 ( .INP(n902), .ZN(n681) );
  INVX0 U1019 ( .INP(n681), .ZN(n682) );
  AND2X1 U1020 ( .IN1(n736), .IN2(n676), .Q(n796) );
  OAI21X1 U1021 ( .IN1(n884), .IN2(n856), .IN3(n519), .QN(g6114) );
  INVX0 U1022 ( .INP(g310), .ZN(n683) );
  INVX0 U1023 ( .INP(n683), .ZN(n684) );
  NBUFFX2 U1024 ( .INP(n919), .Z(n685) );
  NBUFFX2 U1025 ( .INP(n455), .Z(n1014) );
  INVX0 U1026 ( .INP(n773), .ZN(n505) );
  AND2X1 U1027 ( .IN1(n573), .IN2(n182), .Q(n580) );
  NBUFFX2 U1028 ( .INP(g98), .Z(n686) );
  INVX0 U1029 ( .INP(g102), .ZN(n887) );
  OAI221X1 U1030 ( .IN1(n517), .IN2(n505), .IN3(n951), .IN4(g175), .IN5(n970), 
        .QN(n920) );
  INVX0 U1031 ( .INP(g314), .ZN(n687) );
  INVX0 U1032 ( .INP(n687), .ZN(n688) );
  NAND3X1 U1033 ( .IN1(n712), .IN2(n174), .IN3(g684), .QN(n172) );
  XNOR3X1 U1034 ( .IN1(n689), .IN2(n690), .IN3(n792), .Q(n585) );
  XOR2X1 U1035 ( .IN1(g18), .IN2(g14), .Q(n689) );
  XNOR2X1 U1036 ( .IN1(g10), .IN2(g1), .Q(n690) );
  XOR2X2 U1037 ( .IN1(n327), .IN2(g478), .Q(n310) );
  NOR2X0 U1038 ( .IN1(n775), .IN2(n776), .QN(n700) );
  INVX0 U1039 ( .INP(n421), .ZN(n691) );
  NAND2X1 U1040 ( .IN1(n751), .IN2(g79), .QN(n692) );
  NAND2X0 U1041 ( .IN1(n415), .IN2(n691), .QN(n693) );
  AO22X2 U1042 ( .IN1(n21), .IN2(n981), .IN3(n990), .IN4(n708), .Q(g6287) );
  AO22X2 U1043 ( .IN1(n953), .IN2(n1016), .IN3(n564), .IN4(n990), .Q(g5626) );
  AO22X2 U1044 ( .IN1(g694), .IN2(n1016), .IN3(n990), .IN4(n576), .Q(g5533) );
  DELLN1X2 U1045 ( .INP(g41), .Z(n694) );
  INVX0 U1046 ( .INP(n137), .ZN(n695) );
  INVX0 U1047 ( .INP(g59), .ZN(n137) );
  INVX0 U1048 ( .INP(g319), .ZN(n696) );
  DELLN1X2 U1049 ( .INP(g89), .Z(n697) );
  NAND3X0 U1050 ( .IN1(n678), .IN2(n307), .IN3(g282), .QN(n306) );
  AND2X1 U1051 ( .IN1(n264), .IN2(n711), .Q(n175) );
  AND4X1 U1052 ( .IN1(g699), .IN2(n785), .IN3(g702), .IN4(n155), .Q(n264) );
  OAI21X1 U1053 ( .IN1(n781), .IN2(g107), .IN3(n165), .QN(n773) );
  NOR2X0 U1054 ( .IN1(n667), .IN2(n415), .QN(n409) );
  NOR2X0 U1055 ( .IN1(n776), .IN2(n775), .QN(n466) );
  NAND3X1 U1056 ( .IN1(n892), .IN2(n213), .IN3(g694), .QN(n212) );
  INVX0 U1057 ( .INP(g606), .ZN(n701) );
  INVX0 U1058 ( .INP(n701), .ZN(n702) );
  NAND2X0 U1059 ( .IN1(n534), .IN2(n671), .QN(n522) );
  NBUFFX2 U1060 ( .INP(n147), .Z(n703) );
  NBUFFX2 U1061 ( .INP(n165), .Z(n867) );
  NBUFFX2 U1062 ( .INP(g345), .Z(n704) );
  OA22X1 U1063 ( .IN1(g697), .IN2(n762), .IN3(g696), .IN4(n64), .Q(n336) );
  NAND3X1 U1064 ( .IN1(n64), .IN2(n17), .IN3(n803), .QN(n334) );
  OA222X1 U1065 ( .IN1(n713), .IN2(n130), .IN3(n695), .IN4(n420), .IN5(n137), 
        .IN6(n422), .Q(n431) );
  NOR2X0 U1066 ( .IN1(n421), .IN2(n752), .QN(n414) );
  NOR2X0 U1067 ( .IN1(n868), .IN2(g357), .QN(n1015) );
  AO21X1 U1068 ( .IN1(n450), .IN2(n451), .IN3(n6), .Q(n449) );
  AND3X1 U1069 ( .IN1(n265), .IN2(n402), .IN3(n1027), .Q(n705) );
  AND2X1 U1070 ( .IN1(n785), .IN2(n705), .Q(n390) );
  AND2X1 U1071 ( .IN1(g699), .IN2(g702), .Q(n402) );
  OAI21X1 U1072 ( .IN1(n454), .IN2(n460), .IN3(n235), .QN(n864) );
  NAND2X1 U1073 ( .IN1(n828), .IN2(n829), .QN(n561) );
  NBUFFX2 U1074 ( .INP(g338), .Z(n706) );
  NAND3X4 U1075 ( .IN1(n887), .IN2(n541), .IN3(n160), .QN(n182) );
  OR2X1 U1076 ( .IN1(n889), .IN2(n885), .Q(n517) );
  OA22X1 U1077 ( .IN1(g170), .IN2(n885), .IN3(n889), .IN4(n109), .Q(n512) );
  NAND2X0 U1078 ( .IN1(n592), .IN2(g323), .QN(n591) );
  XOR2X1 U1079 ( .IN1(n430), .IN2(g64), .Q(n429) );
  AO21X1 U1080 ( .IN1(n444), .IN2(n445), .IN3(n6), .Q(n443) );
  NAND2X1 U1081 ( .IN1(n1015), .IN2(n464), .QN(n454) );
  NBUFFX2 U1082 ( .INP(n854), .Z(n707) );
  AND2X1 U1083 ( .IN1(n819), .IN2(n138), .Q(n546) );
  NBUFFX2 U1084 ( .INP(n475), .Z(n708) );
  NBUFFX2 U1085 ( .INP(n394), .Z(n991) );
  NOR3X0 U1086 ( .IN1(n463), .IN2(n55), .IN3(n132), .QN(n751) );
  NAND3X1 U1087 ( .IN1(n147), .IN2(n790), .IN3(n1014), .QN(n235) );
  NAND2X0 U1088 ( .IN1(n609), .IN2(n738), .QN(n709) );
  NOR3X0 U1089 ( .IN1(n740), .IN2(n799), .IN3(n476), .QN(g6295) );
  INVX0 U1090 ( .INP(g679), .ZN(n710) );
  INVX0 U1091 ( .INP(g658), .ZN(n120) );
  NBUFFX2 U1092 ( .INP(n265), .Z(n711) );
  OAI221X1 U1093 ( .IN1(g394), .IN2(n713), .IN3(n407), .IN4(n412), .IN5(n919), 
        .QN(n928) );
  NBUFFX2 U1094 ( .INP(n390), .Z(n712) );
  AO21X1 U1095 ( .IN1(n241), .IN2(n696), .IN3(n709), .Q(n713) );
  DELLN2X2 U1096 ( .INP(n609), .Z(n714) );
  NOR2X0 U1097 ( .IN1(g59), .IN2(n665), .QN(n423) );
  NBUFFX2 U1098 ( .INP(n976), .Z(n716) );
  NAND3X0 U1099 ( .IN1(n912), .IN2(n100), .IN3(n1029), .QN(n363) );
  NOR2X0 U1100 ( .IN1(n718), .IN2(n821), .QN(n717) );
  INVX0 U1101 ( .INP(n977), .ZN(n979) );
  IBUFFX16 U1102 ( .INP(n1022), .ZN(n1023) );
  AND3X1 U1103 ( .IN1(n263), .IN2(g687), .IN3(n742), .Q(n847) );
  XOR2X1 U1104 ( .IN1(n418), .IN2(g74), .Q(n417) );
  AND3X1 U1105 ( .IN1(n86), .IN2(g683), .IN3(n397), .Q(n396) );
  NAND3X0 U1106 ( .IN1(n437), .IN2(n436), .IN3(n442), .QN(n441) );
  NBUFFX2 U1107 ( .INP(g642), .Z(n720) );
  NAND2X0 U1108 ( .IN1(n439), .IN2(n443), .QN(g6444) );
  NAND2X0 U1109 ( .IN1(n439), .IN2(n449), .QN(g6440) );
  DELLN2X2 U1110 ( .INP(n868), .Z(n722) );
  OR2X1 U1111 ( .IN1(g338), .IN2(g341), .Q(n723) );
  INVX0 U1112 ( .INP(g40), .ZN(n724) );
  INVX0 U1113 ( .INP(n724), .ZN(g4105) );
  INVX0 U1114 ( .INP(g39), .ZN(n726) );
  INVX0 U1115 ( .INP(n726), .ZN(g4103) );
  INVX0 U1116 ( .INP(g38), .ZN(n728) );
  INVX0 U1117 ( .INP(n728), .ZN(g4102) );
  INVX0 U1118 ( .INP(g37), .ZN(n730) );
  INVX0 U1119 ( .INP(n730), .ZN(g4101) );
  INVX0 U1120 ( .INP(g36), .ZN(n732) );
  INVX0 U1121 ( .INP(n732), .ZN(g4100) );
  INVX0 U1122 ( .INP(g32), .ZN(n734) );
  INVX0 U1123 ( .INP(n734), .ZN(g4099) );
  INVX0 U1124 ( .INP(g314), .ZN(n913) );
  AO21X1 U1125 ( .IN1(n241), .IN2(n696), .IN3(n709), .Q(n854) );
  INVX0 U1126 ( .INP(n534), .ZN(n736) );
  AND4X1 U1127 ( .IN1(n401), .IN2(g675), .IN3(n694), .IN4(n144), .Q(n488) );
  NAND3X0 U1128 ( .IN1(n737), .IN2(n144), .IN3(g675), .QN(g6282) );
  NOR2X0 U1129 ( .IN1(g353), .IN2(g357), .QN(n738) );
  INVX0 U1130 ( .INP(n17), .ZN(n739) );
  NAND2X0 U1131 ( .IN1(n783), .IN2(n827), .QN(n836) );
  AO21X1 U1132 ( .IN1(n700), .IN2(g594), .IN3(n159), .Q(n740) );
  NBUFFX2 U1133 ( .INP(n1024), .Z(n741) );
  NBUFFX2 U1134 ( .INP(n390), .Z(n742) );
  NAND3X1 U1135 ( .IN1(n420), .IN2(n422), .IN3(n435), .QN(n434) );
  NAND2X0 U1136 ( .IN1(n314), .IN2(n317), .QN(n743) );
  AO22X1 U1137 ( .IN1(g642), .IN2(n968), .IN3(g230), .IN4(n880), .Q(n252) );
  DELLN2X2 U1138 ( .INP(n585), .Z(n744) );
  INVX0 U1139 ( .INP(n392), .ZN(n850) );
  NAND2X0 U1140 ( .IN1(n542), .IN2(n921), .QN(n745) );
  NAND2X1 U1141 ( .IN1(n888), .IN2(n794), .QN(n746) );
  NAND2X1 U1142 ( .IN1(n745), .IN2(n746), .QN(n534) );
  NBUFFX2 U1143 ( .INP(n145), .Z(n749) );
  NBUFFX2 U1144 ( .INP(n202), .Z(n843) );
  NBUFFX2 U1145 ( .INP(n172), .Z(n750) );
  NBUFFX2 U1146 ( .INP(n910), .Z(n866) );
  INVX0 U1147 ( .INP(n1024), .ZN(n753) );
  INVX0 U1148 ( .INP(n119), .ZN(n754) );
  INVX0 U1149 ( .INP(n793), .ZN(n755) );
  NBUFFX2 U1150 ( .INP(n57), .Z(n793) );
  NAND2X0 U1151 ( .IN1(n316), .IN2(n320), .QN(n315) );
  NBUFFX2 U1152 ( .INP(n686), .Z(n757) );
  INVX0 U1153 ( .INP(n977), .ZN(n978) );
  INVX0 U1154 ( .INP(g345), .ZN(n103) );
  NAND2X0 U1155 ( .IN1(g161), .IN2(n796), .QN(n758) );
  NAND2X0 U1156 ( .IN1(n796), .IN2(g161), .QN(n509) );
  AO221X1 U1157 ( .IN1(n313), .IN2(n852), .IN3(n314), .IN4(g211), .IN5(n15), 
        .Q(n759) );
  NBUFFX2 U1158 ( .INP(n119), .Z(n760) );
  NBUFFX2 U1159 ( .INP(n364), .Z(n761) );
  DELLN1X2 U1160 ( .INP(g276), .Z(n762) );
  NBUFFX2 U1161 ( .INP(n631), .Z(n763) );
  NBUFFX2 U1162 ( .INP(n958), .Z(n764) );
  AND2X1 U1163 ( .IN1(n334), .IN2(n34), .Q(n765) );
  INVX0 U1164 ( .INP(g638), .ZN(n766) );
  NBUFFX2 U1165 ( .INP(n786), .Z(n767) );
  INVX0 U1166 ( .INP(n363), .ZN(n768) );
  INVX0 U1167 ( .INP(n768), .ZN(n769) );
  AO22X2 U1168 ( .IN1(n981), .IN2(n1010), .IN3(n563), .IN4(n64), .Q(g5532) );
  NAND2X1 U1169 ( .IN1(n194), .IN2(n666), .QN(n180) );
  AOI222X1 U1170 ( .IN1(n862), .IN2(n196), .IN3(n197), .IN4(n880), .IN5(n2), 
        .IN6(n52), .QN(n170) );
  NBUFFX2 U1171 ( .INP(n369), .Z(n770) );
  NAND2X1 U1172 ( .IN1(n373), .IN2(n717), .QN(g6480) );
  NAND2X1 U1173 ( .IN1(n237), .IN2(n670), .QN(n236) );
  NAND3X0 U1174 ( .IN1(n886), .IN2(n128), .IN3(g682), .QN(n379) );
  AO22X1 U1175 ( .IN1(g697), .IN2(n1039), .IN3(n179), .IN4(g269), .Q(g6794) );
  AO22X1 U1176 ( .IN1(n855), .IN2(g434), .IN3(n865), .IN4(g430), .Q(n288) );
  INVX0 U1177 ( .INP(n1041), .ZN(n772) );
  NBUFFX2 U1178 ( .INP(n179), .Z(n903) );
  AO22X1 U1179 ( .IN1(n855), .IN2(g441), .IN3(n971), .IN4(g422), .Q(n353) );
  AO22X1 U1180 ( .IN1(n764), .IN2(g445), .IN3(n971), .IN4(g418), .Q(n357) );
  AO22X1 U1181 ( .IN1(n764), .IN2(g437), .IN3(n971), .IN4(g426), .Q(n295) );
  AND2X4 U1182 ( .IN1(n462), .IN2(n459), .Q(n774) );
  AO21X1 U1183 ( .IN1(n1035), .IN2(n875), .IN3(n863), .Q(n375) );
  NAND2X0 U1184 ( .IN1(n473), .IN2(g586), .QN(n775) );
  OR2X1 U1185 ( .IN1(n777), .IN2(n88), .Q(n776) );
  INVX0 U1186 ( .INP(g590), .ZN(n777) );
  INVX0 U1187 ( .INP(n778), .ZN(n779) );
  AND2X1 U1188 ( .IN1(n864), .IN2(n780), .Q(n791) );
  INVX0 U1189 ( .INP(n791), .ZN(n439) );
  AND3X1 U1190 ( .IN1(n143), .IN2(n160), .IN3(n541), .Q(n781) );
  OR2X1 U1191 ( .IN1(n548), .IN2(n540), .Q(n783) );
  AO22X1 U1192 ( .IN1(n881), .IN2(n739), .IN3(g520), .IN4(n716), .Q(g6309) );
  AO21X1 U1193 ( .IN1(n529), .IN2(n530), .IN3(n884), .Q(n528) );
  AND3X1 U1194 ( .IN1(n364), .IN2(n362), .IN3(n363), .Q(n784) );
  OAI222X1 U1195 ( .IN1(n362), .IN2(n97), .IN3(n83), .IN4(n769), .IN5(n43), 
        .IN6(n761), .QN(n998) );
  OA222X1 U1196 ( .IN1(n362), .IN2(n99), .IN3(n92), .IN4(n769), .IN5(n47), 
        .IN6(n761), .Q(n367) );
  OA222X1 U1197 ( .IN1(n798), .IN2(n27), .IN3(n1010), .IN4(n363), .IN5(n121), 
        .IN6(n364), .Q(n372) );
  OA21X1 U1198 ( .IN1(n694), .IN2(n586), .IN3(g676), .Q(n785) );
  OA21X1 U1199 ( .IN1(n694), .IN2(n771), .IN3(g676), .Q(n401) );
  NAND3X1 U1200 ( .IN1(n742), .IN2(n793), .IN3(n174), .QN(n202) );
  OA21X1 U1201 ( .IN1(n460), .IN2(n454), .IN3(n235), .Q(n786) );
  NBUFFX2 U1202 ( .INP(g205), .Z(n787) );
  AO22X2 U1203 ( .IN1(g548), .IN2(n301), .IN3(n960), .IN4(n759), .Q(g6788) );
  AND4X1 U1204 ( .IN1(n836), .IN2(n680), .IN3(n543), .IN4(n827), .Q(n902) );
  OR2X1 U1205 ( .IN1(n152), .IN2(g310), .Q(n788) );
  NBUFFX2 U1206 ( .INP(n631), .Z(n1033) );
  NBUFFX2 U1207 ( .INP(n631), .Z(n1034) );
  AO22X2 U1208 ( .IN1(g696), .IN2(n1017), .IN3(n990), .IN4(n743), .Q(g6791) );
  AND2X1 U1209 ( .IN1(n822), .IN2(n12), .Q(n571) );
  XNOR3X1 U1210 ( .IN1(g24), .IN2(g2), .IN3(n830), .Q(n792) );
  XOR2X1 U1211 ( .IN1(g6), .IN2(g28), .Q(n830) );
  AO21X1 U1212 ( .IN1(n59), .IN2(n849), .IN3(n809), .Q(n577) );
  NBUFFX2 U1213 ( .INP(n459), .Z(n810) );
  DELLN1X2 U1214 ( .INP(g94), .Z(n794) );
  NBUFFX2 U1215 ( .INP(n534), .Z(n795) );
  OR3X1 U1216 ( .IN1(n106), .IN2(n795), .IN3(n133), .Q(n523) );
  INVX0 U1217 ( .INP(n362), .ZN(n797) );
  INVX0 U1218 ( .INP(n797), .ZN(n798) );
  NAND2X1 U1219 ( .IN1(n681), .IN2(n528), .QN(g6109) );
  NAND3X1 U1220 ( .IN1(n531), .IN2(n969), .IN3(n532), .QN(n530) );
  OA222X1 U1221 ( .IN1(n135), .IN2(n798), .IN3(n1016), .IN4(n769), .IN5(n102), 
        .IN6(n761), .Q(n382) );
  AND2X1 U1222 ( .IN1(n29), .IN2(n800), .Q(g6299) );
  OR2X1 U1223 ( .IN1(n799), .IN2(g586), .Q(n472) );
  NBUFFX2 U1224 ( .INP(g277), .Z(n803) );
  INVX0 U1225 ( .INP(g306), .ZN(n804) );
  INVX0 U1226 ( .INP(n804), .ZN(n805) );
  NBUFFX2 U1227 ( .INP(n339), .Z(n806) );
  INVX0 U1228 ( .INP(n573), .ZN(n807) );
  NAND3X0 U1229 ( .IN1(n383), .IN2(n668), .IN3(n380), .QN(g6479) );
  INVX0 U1230 ( .INP(n808), .ZN(n809) );
  INVX0 U1231 ( .INP(n458), .ZN(n811) );
  NOR2X0 U1232 ( .IN1(n984), .IN2(n964), .QN(n813) );
  AND2X1 U1233 ( .IN1(n813), .IN2(n814), .Q(n645) );
  NOR2X0 U1234 ( .IN1(n548), .IN2(n540), .QN(n819) );
  NAND2X1 U1235 ( .IN1(n372), .IN2(n371), .QN(n821) );
  NOR2X0 U1236 ( .IN1(n566), .IN2(n1016), .QN(n822) );
  NOR2X0 U1237 ( .IN1(n568), .IN2(n669), .QN(n480) );
  DELLN2X2 U1238 ( .INP(g28), .Z(n825) );
  INVX0 U1239 ( .INP(n333), .ZN(n828) );
  NBUFFX2 U1240 ( .INP(n299), .Z(n826) );
  AND2X1 U1241 ( .IN1(g278), .IN2(g279), .Q(n829) );
  INVX0 U1242 ( .INP(n686), .ZN(n831) );
  INVX0 U1243 ( .INP(n831), .ZN(n832) );
  AND2X1 U1244 ( .IN1(n311), .IN2(g282), .Q(n833) );
  AND2X1 U1245 ( .IN1(n310), .IN2(n833), .Q(n305) );
  AO22X2 U1246 ( .IN1(g551), .IN2(n301), .IN3(n960), .IN4(n178), .Q(g6789) );
  AO22X2 U1247 ( .IN1(n846), .IN2(n1011), .IN3(n992), .IN4(n178), .Q(g6793) );
  NAND2X1 U1248 ( .IN1(n303), .IN2(n306), .QN(n178) );
  DELLN2X2 U1249 ( .INP(n621), .Z(n834) );
  AO22X1 U1250 ( .IN1(n1040), .IN2(n755), .IN3(n772), .IN4(n279), .Q(n282) );
  NBUFFX2 U1251 ( .INP(g699), .Z(g1293) );
  INVX0 U1252 ( .INP(n860), .ZN(n857) );
  AND4X1 U1253 ( .IN1(n633), .IN2(n634), .IN3(n635), .IN4(n636), .Q(n837) );
  INVX0 U1254 ( .INP(n927), .ZN(n961) );
  INVX0 U1255 ( .INP(g694), .ZN(n841) );
  INVX0 U1256 ( .INP(n841), .ZN(n842) );
  NBUFFX2 U1257 ( .INP(n326), .Z(n844) );
  NOR2X0 U1258 ( .IN1(n311), .IN2(n481), .QN(n326) );
  INVX0 U1259 ( .INP(n747), .ZN(n845) );
  NAND2X1 U1260 ( .IN1(n899), .IN2(n672), .QN(g6937) );
  NBUFFX2 U1261 ( .INP(g696), .Z(n846) );
  NAND2X1 U1262 ( .IN1(g123), .IN2(n166), .QN(n901) );
  AND2X1 U1263 ( .IN1(g578), .IN2(n878), .Q(n848) );
  NOR3X0 U1264 ( .IN1(n561), .IN2(g280), .IN3(n77), .QN(n481) );
  INVX0 U1265 ( .INP(n850), .ZN(n851) );
  AND4X1 U1266 ( .IN1(n770), .IN2(n387), .IN3(n378), .IN4(n376), .Q(n853) );
  NAND3X1 U1267 ( .IN1(g301), .IN2(n154), .IN3(n688), .QN(n456) );
  NBUFFX2 U1268 ( .INP(n958), .Z(n855) );
  AND2X1 U1269 ( .IN1(n454), .IN2(n1013), .Q(n896) );
  XNOR2X1 U1270 ( .IN1(n109), .IN2(n920), .Q(n856) );
  DELLN1X2 U1271 ( .INP(n408), .Z(n869) );
  AOI21X1 U1272 ( .IN1(n536), .IN2(n537), .IN3(n845), .QN(n858) );
  AND2X1 U1273 ( .IN1(n872), .IN2(n103), .Q(n589) );
  XNOR2X1 U1274 ( .IN1(g84), .IN2(n1028), .Q(n859) );
  NBUFFX2 U1275 ( .INP(n24), .Z(n861) );
  NBUFFX2 U1276 ( .INP(n1031), .Z(n862) );
  INVX0 U1277 ( .INP(n284), .ZN(n863) );
  INVX0 U1278 ( .INP(g658), .ZN(n1038) );
  AO22X1 U1279 ( .IN1(n892), .IN2(n1031), .IN3(g224), .IN4(n880), .Q(n256) );
  INVX0 U1280 ( .INP(n439), .ZN(n1025) );
  NAND3X1 U1281 ( .IN1(n760), .IN2(n136), .IN3(g205), .QN(n345) );
  NBUFFX2 U1282 ( .INP(n972), .Z(n865) );
  INVX0 U1283 ( .INP(n715), .ZN(n972) );
  AO22X1 U1284 ( .IN1(g650), .IN2(n1031), .IN3(g248), .IN4(n879), .Q(n279) );
  NAND2X0 U1285 ( .IN1(n609), .IN2(n101), .QN(n868) );
  OA222X2 U1286 ( .IN1(n1012), .IN2(n62), .IN3(n80), .IN4(n420), .IN5(n421), 
        .IN6(n422), .Q(n419) );
  INVX0 U1287 ( .INP(g639), .ZN(n870) );
  NOR2X0 U1288 ( .IN1(n140), .IN2(n867), .QN(n166) );
  NAND2X0 U1289 ( .IN1(n164), .IN2(n867), .QN(n900) );
  XNOR2X1 U1290 ( .IN1(n511), .IN2(g179), .Q(n871) );
  AO22X1 U1291 ( .IN1(n688), .IN2(n805), .IN3(n788), .IN4(n913), .Q(n462) );
  NOR2X0 U1292 ( .IN1(n723), .IN2(g349), .QN(n872) );
  NAND2X0 U1293 ( .IN1(n64), .IN2(n803), .QN(n873) );
  NAND2X0 U1294 ( .IN1(n136), .IN2(n874), .QN(n332) );
  INVX0 U1295 ( .INP(n873), .ZN(n874) );
  NBUFFX2 U1296 ( .INP(g691), .Z(n875) );
  NAND2X1 U1297 ( .IN1(n328), .IN2(n329), .QN(n327) );
  NOR3X0 U1298 ( .IN1(n621), .IN2(g139), .IN3(g135), .QN(n165) );
  AND2X1 U1299 ( .IN1(n624), .IN2(g625), .Q(n877) );
  AND2X1 U1300 ( .IN1(g631), .IN2(g628), .Q(n878) );
  INVX0 U1301 ( .INP(n1037), .ZN(n879) );
  INVX0 U1302 ( .INP(n976), .ZN(n881) );
  INVX0 U1303 ( .INP(n976), .ZN(n882) );
  INVX0 U1304 ( .INP(n469), .ZN(n883) );
  NAND2X0 U1305 ( .IN1(g639), .IN2(n649), .QN(g3828) );
  AO21X1 U1306 ( .IN1(n777), .IN2(n883), .IN3(n922), .Q(n465) );
  INVX0 U1307 ( .INP(n747), .ZN(n884) );
  NOR2X0 U1308 ( .IN1(n820), .IN2(g161), .QN(n885) );
  NOR2X0 U1309 ( .IN1(n522), .IN2(g161), .QN(n513) );
  XNOR2X2 U1310 ( .IN1(n585), .IN2(g48), .Q(n586) );
  INVX0 U1311 ( .INP(n887), .ZN(n888) );
  NOR2X0 U1312 ( .IN1(n134), .IN2(n523), .QN(n889) );
  INVX0 U1313 ( .INP(n519), .ZN(n890) );
  INVX0 U1314 ( .INP(n902), .ZN(n519) );
  INVX0 U1315 ( .INP(g634), .ZN(n891) );
  NOR2X0 U1316 ( .IN1(n923), .IN2(n904), .QN(n630) );
  NAND2X1 U1317 ( .IN1(n967), .IN2(g662), .QN(n171) );
  NBUFFX2 U1318 ( .INP(n896), .Z(n894) );
  OAI21X1 U1319 ( .IN1(n452), .IN2(n894), .IN3(g361), .QN(n450) );
  INVX0 U1320 ( .INP(n474), .ZN(n895) );
  AO21X1 U1321 ( .IN1(n88), .IN2(n779), .IN3(n469), .Q(n467) );
  AO21X1 U1322 ( .IN1(n105), .IN2(n650), .IN3(n651), .Q(n649) );
  AO22X1 U1323 ( .IN1(g554), .IN2(n301), .IN3(n960), .IN4(n903), .Q(g6790) );
  INVX0 U1324 ( .INP(g697), .ZN(n897) );
  INVX0 U1325 ( .INP(n897), .ZN(n898) );
  NAND2X1 U1326 ( .IN1(n140), .IN2(n163), .QN(n899) );
  NAND2X1 U1327 ( .IN1(n335), .IN2(n765), .QN(n328) );
  XNOR2X2 U1328 ( .IN1(g6794), .IN2(n926), .Q(n237) );
  NAND2X0 U1329 ( .IN1(n286), .IN2(n673), .QN(g6845) );
  NOR2X0 U1330 ( .IN1(n923), .IN2(n924), .QN(n647) );
  INVX0 U1331 ( .INP(g619), .ZN(n905) );
  NAND3X0 U1332 ( .IN1(n161), .IN2(n141), .IN3(n832), .QN(n193) );
  INVX0 U1333 ( .INP(g205), .ZN(n906) );
  OR2X1 U1334 ( .IN1(n924), .IN2(n905), .Q(n904) );
  OR2X1 U1335 ( .IN1(n75), .IN2(n907), .Q(n908) );
  INVX0 U1336 ( .INP(g204), .ZN(n907) );
  OR2X1 U1337 ( .IN1(n906), .IN2(n907), .Q(n346) );
  INVX0 U1338 ( .INP(n12), .ZN(n909) );
  NAND2X0 U1339 ( .IN1(n853), .IN2(n385), .QN(n910) );
  INVX0 U1340 ( .INP(n911), .ZN(n912) );
  INVX0 U1341 ( .INP(n984), .ZN(n986) );
  INVX0 U1342 ( .INP(n964), .ZN(n966) );
  NBUFFX2 U1343 ( .INP(n550), .Z(n914) );
  NBUFFX2 U1344 ( .INP(n550), .Z(n915) );
  NBUFFX2 U1345 ( .INP(n550), .Z(n916) );
  NBUFFX2 U1346 ( .INP(n854), .Z(n1013) );
  NBUFFX2 U1347 ( .INP(n141), .Z(n921) );
  INVX0 U1348 ( .INP(n31), .ZN(n918) );
  NAND2X0 U1349 ( .IN1(n454), .IN2(n707), .QN(n919) );
  NAND3X1 U1350 ( .IN1(n742), .IN2(n91), .IN3(g689), .QN(n389) );
  NAND2X0 U1351 ( .IN1(g602), .IN2(g610), .QN(n923) );
  INVX0 U1352 ( .INP(g616), .ZN(n925) );
  INVX0 U1353 ( .INP(n299), .ZN(n68) );
  INVX0 U1354 ( .INP(n1022), .ZN(n1024) );
  NBUFFX2 U1355 ( .INP(n123), .Z(n1017) );
  NBUFFX2 U1356 ( .INP(n123), .Z(n1016) );
  NOR3X0 U1357 ( .IN1(n1041), .IN2(n918), .IN3(n559), .QN(n563) );
  INVX0 U1358 ( .INP(n566), .ZN(n13) );
  INVX0 U1359 ( .INP(n559), .ZN(n32) );
  INVX0 U1360 ( .INP(n323), .ZN(n12) );
  INVX0 U1361 ( .INP(n312), .ZN(n31) );
  NBUFFX2 U1362 ( .INP(n763), .Z(n1032) );
  INVX0 U1363 ( .INP(n166), .ZN(n35) );
  NOR2X0 U1364 ( .IN1(n42), .IN2(n158), .QN(n219) );
  INVX0 U1365 ( .INP(n956), .ZN(n958) );
  NBUFFX2 U1366 ( .INP(n488), .Z(n1045) );
  INVX0 U1367 ( .INP(n471), .ZN(n20) );
  NBUFFX2 U1368 ( .INP(n488), .Z(n1046) );
  NBUFFX2 U1369 ( .INP(n488), .Z(n1044) );
  INVX0 U1370 ( .INP(n475), .ZN(n21) );
  INVX0 U1371 ( .INP(n545), .ZN(n987) );
  NOR2X0 U1372 ( .IN1(n986), .IN2(n966), .QN(n213) );
  INVX0 U1373 ( .INP(n578), .ZN(n74) );
  INVX0 U1374 ( .INP(n579), .ZN(n82) );
  NAND2X0 U1375 ( .IN1(n860), .IN2(n305), .QN(n304) );
  NAND2X0 U1376 ( .IN1(n230), .IN2(n231), .QN(n655) );
  INVX0 U1377 ( .INP(n309), .ZN(n33) );
  INVX0 U1378 ( .INP(n320), .ZN(n14) );
  NOR2X0 U1379 ( .IN1(n151), .IN2(n458), .QN(n457) );
  INVX0 U1380 ( .INP(n927), .ZN(n962) );
  INVX0 U1381 ( .INP(n200), .ZN(n52) );
  NAND3X0 U1382 ( .IN1(n99), .IN2(n97), .IN3(n837), .QN(n631) );
  INVX0 U1383 ( .INP(n250), .ZN(n41) );
  INVX0 U1384 ( .INP(n369), .ZN(n24) );
  INVX0 U1385 ( .INP(n545), .ZN(n69) );
  INVX0 U1386 ( .INP(n985), .ZN(n158) );
  OA21X1 U1387 ( .IN1(n607), .IN2(n67), .IN3(n826), .Q(g5050) );
  NOR2X0 U1388 ( .IN1(n714), .IN2(n101), .QN(n607) );
  INVX0 U1389 ( .INP(g598), .ZN(n42) );
  INVX0 U1390 ( .INP(n773), .ZN(n949) );
  INVX0 U1391 ( .INP(n252), .ZN(n112) );
  INVX0 U1392 ( .INP(n538), .ZN(n37) );
  INVX0 U1393 ( .INP(n531), .ZN(n38) );
  NAND2X0 U1394 ( .IN1(n1044), .IN2(n49), .QN(g6110) );
  INVX0 U1395 ( .INP(g6658), .ZN(n49) );
  NAND3X0 U1396 ( .IN1(g693), .IN2(n76), .IN3(n219), .QN(n215) );
  NOR2X0 U1397 ( .IN1(n214), .IN2(n653), .QN(g3454) );
  INVX0 U1398 ( .INP(n930), .ZN(n976) );
  AND4X1 U1399 ( .IN1(n244), .IN2(n811), .IN3(n810), .IN4(n242), .Q(n300) );
  NAND2X0 U1400 ( .IN1(n71), .IN2(n625), .QN(g4607) );
  NAND2X0 U1401 ( .IN1(n124), .IN2(n628), .QN(g4497) );
  INVX0 U1402 ( .INP(n810), .ZN(n151) );
  INVX0 U1403 ( .INP(n186), .ZN(g1802) );
  NAND2X0 U1404 ( .IN1(n263), .IN2(n175), .QN(n261) );
  INVX0 U1405 ( .INP(n311), .ZN(n78) );
  INVX0 U1406 ( .INP(n322), .ZN(n58) );
  INVX0 U1407 ( .INP(n498), .ZN(n115) );
  INVX0 U1408 ( .INP(n239), .ZN(n148) );
  INVX0 U1409 ( .INP(n952), .ZN(n953) );
  INVX0 U1410 ( .INP(n954), .ZN(n955) );
  INVX0 U1411 ( .INP(n162), .ZN(n23) );
  INVX0 U1412 ( .INP(n964), .ZN(n965) );
  INVX0 U1413 ( .INP(n596), .ZN(n66) );
  INVX0 U1414 ( .INP(g281), .ZN(n77) );
  INVX0 U1415 ( .INP(g188), .ZN(n51) );
  INVX0 U1416 ( .INP(g698), .ZN(n91) );
  OA22X1 U1417 ( .IN1(g332), .IN2(n240), .IN3(n242), .IN4(n8), .Q(n926) );
  INVX0 U1418 ( .INP(g161), .ZN(n134) );
  NOR2X0 U1419 ( .IN1(n316), .IN2(n117), .QN(n313) );
  INVX0 U1420 ( .INP(n315), .ZN(n15) );
  INVX0 U1421 ( .INP(g210), .ZN(n117) );
  INVX0 U1422 ( .INP(g179), .ZN(n45) );
  NOR2X0 U1423 ( .IN1(n305), .IN2(n73), .QN(n302) );
  INVX0 U1424 ( .INP(n304), .ZN(n16) );
  INVX0 U1425 ( .INP(g282), .ZN(n73) );
  NAND2X0 U1426 ( .IN1(g281), .IN2(n553), .QN(n309) );
  NAND2X0 U1427 ( .IN1(g209), .IN2(n556), .QN(n320) );
  NOR2X0 U1428 ( .IN1(g123), .IN2(n167), .QN(n164) );
  OA21X1 U1429 ( .IN1(n787), .IN2(n754), .IN3(n346), .Q(n572) );
  NAND2X1 U1430 ( .IN1(n53), .IN2(g54), .QN(n422) );
  INVX0 U1431 ( .INP(n436), .ZN(n53) );
  NOR2X0 U1432 ( .IN1(n757), .IN2(g94), .QN(n541) );
  OA222X1 U1433 ( .IN1(n1012), .IN2(n95), .IN3(n420), .IN4(n427), .IN5(n422), 
        .IN6(n428), .Q(n426) );
  AO21X1 U1434 ( .IN1(n756), .IN2(n981), .IN3(n863), .Q(n384) );
  NOR2X0 U1435 ( .IN1(g654), .IN2(n611), .QN(n610) );
  NOR2X0 U1436 ( .IN1(n616), .IN2(g650), .QN(n615) );
  NAND2X0 U1437 ( .IN1(n739), .IN2(n756), .QN(n350) );
  NAND2X0 U1438 ( .IN1(n846), .IN2(n756), .QN(n292) );
  NAND2X0 U1439 ( .IN1(n842), .IN2(n1035), .QN(n354) );
  INVX0 U1440 ( .INP(g337), .ZN(n1005) );
  NOR2X0 U1441 ( .IN1(n991), .IN2(n395), .QN(n393) );
  INVX0 U1442 ( .INP(g691), .ZN(n136) );
  NAND2X0 U1443 ( .IN1(n314), .IN2(n317), .QN(n230) );
  NAND2X0 U1444 ( .IN1(n319), .IN2(n58), .QN(n318) );
  INVX0 U1445 ( .INP(n198), .ZN(n2) );
  OA21X1 U1446 ( .IN1(n803), .IN2(n762), .IN3(n917), .Q(n569) );
  NOR2X0 U1447 ( .IN1(n555), .IN2(n1009), .QN(n554) );
  INVX0 U1448 ( .INP(g353), .ZN(n101) );
  NAND2X1 U1449 ( .IN1(n341), .IN2(n342), .QN(n340) );
  OR2X1 U1450 ( .IN1(n1012), .IN2(g366), .Q(n453) );
  NAND2X0 U1451 ( .IN1(n308), .IN2(n78), .QN(n307) );
  XNOR2X1 U1452 ( .IN1(g79), .IN2(n928), .Q(n410) );
  XOR2X1 U1453 ( .IN1(g54), .IN2(n929), .Q(n438) );
  OA21X1 U1454 ( .IN1(n558), .IN2(n559), .IN3(n31), .Q(n557) );
  OA21X1 U1455 ( .IN1(n565), .IN2(n566), .IN3(n12), .Q(n564) );
  AOI22X1 U1456 ( .IN1(g680), .IN2(n1036), .IN3(n989), .IN4(n256), .QN(n271)
         );
  INVX0 U1457 ( .INP(g89), .ZN(n160) );
  NAND2X0 U1458 ( .IN1(g361), .IN2(n453), .QN(n452) );
  NOR4X0 U1459 ( .IN1(n637), .IN2(n638), .IN3(n639), .IN4(n640), .QN(n636) );
  INVX0 U1460 ( .INP(g301), .ZN(n147) );
  INVX0 U1461 ( .INP(g94), .ZN(n161) );
  INVX0 U1462 ( .INP(g319), .ZN(n154) );
  INVX0 U1463 ( .INP(g6690), .ZN(n79) );
  NOR2X0 U1464 ( .IN1(n627), .IN2(g646), .QN(n626) );
  INVX0 U1465 ( .INP(g639), .ZN(n159) );
  NOR2X0 U1466 ( .IN1(g332), .IN2(n300), .QN(n297) );
  INVX0 U1467 ( .INP(n834), .ZN(n40) );
  NAND2X0 U1468 ( .IN1(n587), .IN2(n826), .QN(g5323) );
  NAND2X0 U1469 ( .IN1(n614), .IN2(n166), .QN(g4773) );
  NAND2X0 U1470 ( .IN1(g698), .IN2(g689), .QN(n391) );
  NAND2X0 U1471 ( .IN1(n97), .IN2(n485), .QN(n484) );
  NAND3X0 U1472 ( .IN1(n486), .IN2(n99), .IN3(n960), .QN(n485) );
  NAND2X0 U1473 ( .IN1(g152), .IN2(n532), .QN(n531) );
  AND2X1 U1474 ( .IN1(n487), .IN2(g677), .Q(n930) );
  INVX0 U1475 ( .INP(g135), .ZN(n129) );
  INVX0 U1476 ( .INP(g685), .ZN(n72) );
  NAND2X0 U1477 ( .IN1(g143), .IN2(n539), .QN(n538) );
  INVX0 U1478 ( .INP(g306), .ZN(n152) );
  AOI22X1 U1479 ( .IN1(g678), .IN2(n1036), .IN3(n989), .IN4(n255), .QN(n272)
         );
  NAND2X0 U1480 ( .IN1(g679), .IN2(n198), .QN(n199) );
  AOI222X1 U1481 ( .IN1(n971), .IN2(g410), .IN3(n24), .IN4(g508), .IN5(n855), 
        .IN6(g453), .QN(n366) );
  INVX0 U1482 ( .INP(g6684), .ZN(n118) );
  INVX0 U1483 ( .INP(g6691), .ZN(n127) );
  INVX0 U1484 ( .INP(g6689), .ZN(n50) );
  NOR2X0 U1485 ( .IN1(g74), .IN2(g54), .QN(n461) );
  NOR2X0 U1486 ( .IN1(n702), .IN2(n645), .QN(n644) );
  INVX0 U1487 ( .INP(g638), .ZN(n111) );
  NAND2X0 U1488 ( .IN1(n108), .IN2(n324), .QN(g6704) );
  NAND2X0 U1489 ( .IN1(n1045), .IN2(n90), .QN(g6185) );
  INVX0 U1490 ( .INP(g6685), .ZN(n90) );
  NAND2X0 U1491 ( .IN1(n1046), .IN2(n126), .QN(g6170) );
  INVX0 U1492 ( .INP(g6688), .ZN(n126) );
  NAND2X0 U1493 ( .IN1(n1045), .IN2(n65), .QN(g6167) );
  INVX0 U1494 ( .INP(g6686), .ZN(n65) );
  INVX0 U1495 ( .INP(g679), .ZN(n104) );
  INVX0 U1496 ( .INP(g551), .ZN(n47) );
  INVX0 U1497 ( .INP(g293), .ZN(n92) );
  INVX0 U1498 ( .INP(g204), .ZN(n119) );
  INVX0 U1499 ( .INP(n543), .ZN(n138) );
  INVX0 U1500 ( .INP(g276), .ZN(n64) );
  NOR2X0 U1501 ( .IN1(g681), .IN2(g682), .QN(n398) );
  INVX0 U1502 ( .INP(g695), .ZN(n17) );
  INVX0 U1503 ( .INP(g143), .ZN(n106) );
  NOR2X0 U1504 ( .IN1(n20), .IN2(n479), .QN(n478) );
  INVX0 U1505 ( .INP(g541), .ZN(n97) );
  INVX0 U1506 ( .INP(g682), .ZN(n48) );
  INVX0 U1507 ( .INP(g278), .ZN(n34) );
  NAND2X0 U1508 ( .IN1(n44), .IN2(n337), .QN(g6702) );
  NAND2X0 U1509 ( .IN1(g54), .IN2(g74), .QN(n463) );
  INVX0 U1510 ( .INP(g457), .ZN(n81) );
  INVX0 U1511 ( .INP(g461), .ZN(n18) );
  INVX0 U1512 ( .INP(g634), .ZN(n76) );
  INVX0 U1513 ( .INP(g536), .ZN(n99) );
  INVX0 U1514 ( .INP(g332), .ZN(n8) );
  NOR2X0 U1515 ( .IN1(n214), .IN2(n720), .QN(n648) );
  INVX0 U1516 ( .INP(g683), .ZN(n100) );
  INVX0 U1517 ( .INP(g361), .ZN(n55) );
  NAND2X0 U1518 ( .IN1(g688), .IN2(n26), .QN(n395) );
  INVX0 U1519 ( .INP(n391), .ZN(n26) );
  INVX0 U1520 ( .INP(g280), .ZN(n113) );
  INVX0 U1521 ( .INP(g152), .ZN(n133) );
  INVX0 U1522 ( .INP(g208), .ZN(n59) );
  INVX0 U1523 ( .INP(g206), .ZN(n75) );
  INVX0 U1524 ( .INP(g123), .ZN(n11) );
  NOR2X0 U1525 ( .IN1(g590), .IN2(n89), .QN(n491) );
  NOR3X0 U1526 ( .IN1(n159), .IN2(n647), .IN3(n652), .QN(g3768) );
  NOR3X0 U1527 ( .IN1(n159), .IN2(n604), .IN3(n612), .QN(g4872) );
  NOR3X0 U1528 ( .IN1(n870), .IN2(n613), .IN3(n623), .QN(g4687) );
  NOR3X0 U1529 ( .IN1(n870), .IN2(n674), .IN3(n603), .QN(g5167) );
  INVX0 U1530 ( .INP(g107), .ZN(n143) );
  AO221X1 U1531 ( .IN1(n953), .IN2(n116), .IN3(g578), .IN4(n955), .IN5(g582), 
        .Q(n495) );
  NAND2X1 U1532 ( .IN1(n115), .IN2(n980), .QN(n496) );
  INVX0 U1533 ( .INP(g578), .ZN(n116) );
  NAND2X0 U1534 ( .IN1(g582), .IN2(g578), .QN(n498) );
  INVX0 U1535 ( .INP(g170), .ZN(n109) );
  INVX0 U1536 ( .INP(g678), .ZN(n4) );
  INVX0 U1537 ( .INP(g49), .ZN(n132) );
  INVX0 U1538 ( .INP(g677), .ZN(n128) );
  NAND2X0 U1539 ( .IN1(n688), .IN2(n684), .QN(n244) );
  INVX0 U1540 ( .INP(g687), .ZN(n94) );
  INVX0 U1541 ( .INP(g22), .ZN(n144) );
  DELLN1X2 U1542 ( .INP(g22), .Z(g4104) );
  NAND2X0 U1543 ( .IN1(g638), .IN2(n985), .QN(g3599) );
  INVX0 U1544 ( .INP(g681), .ZN(n63) );
  NOR2X0 U1545 ( .IN1(n228), .IN2(n229), .QN(n226) );
  NAND2X0 U1546 ( .IN1(g64), .IN2(n695), .QN(n428) );
  OR2X1 U1547 ( .IN1(g672), .IN2(n931), .Q(g5231) );
  NOR3X0 U1548 ( .IN1(g22), .IN2(g4110), .IN3(n801), .QN(n931) );
  XOR3X1 U1549 ( .IN1(n932), .IN2(n582), .IN3(n933), .Q(n162) );
  XNOR2X1 U1550 ( .IN1(g48), .IN2(g4105), .Q(n932) );
  INVX0 U1551 ( .INP(g465), .ZN(n27) );
  INVX0 U1552 ( .INP(g6687), .ZN(n84) );
  INVX0 U1553 ( .INP(g574), .ZN(n88) );
  INVX0 U1554 ( .INP(g114), .ZN(n124) );
  INVX0 U1555 ( .INP(g586), .ZN(n89) );
  INVX0 U1556 ( .INP(g492), .ZN(n108) );
  INVX0 U1557 ( .INP(g496), .ZN(n44) );
  INVX0 U1558 ( .INP(g686), .ZN(n110) );
  INVX0 U1559 ( .INP(g386), .ZN(n95) );
  INVX0 U1560 ( .INP(g390), .ZN(n62) );
  INVX0 U1561 ( .INP(g382), .ZN(n130) );
  AND3X1 U1562 ( .IN1(g639), .IN2(n650), .IN3(n654), .Q(g2670) );
  NOR2X0 U1563 ( .IN1(g266), .IN2(n156), .QN(g3910) );
  INVX0 U1564 ( .INP(g45), .ZN(n156) );
  INVX0 U1565 ( .INP(g111), .ZN(n125) );
  INVX0 U1566 ( .INP(g500), .ZN(n122) );
  INVX0 U1567 ( .INP(g504), .ZN(n96) );
  INVX0 U1568 ( .INP(g398), .ZN(n56) );
  INVX0 U1569 ( .INP(g297), .ZN(n83) );
  INVX0 U1570 ( .INP(g554), .ZN(n43) );
  INVX0 U1571 ( .INP(g266), .ZN(n131) );
  INVX0 U1572 ( .INP(g548), .ZN(n121) );
  INVX0 U1573 ( .INP(g545), .ZN(n102) );
  NBUFFX2 U1574 ( .INP(g23), .Z(g4098) );
  DELLN1X2 U1575 ( .INP(g42), .Z(g4106) );
  NBUFFX2 U1576 ( .INP(g44), .Z(g4107) );
  DELLN1X2 U1577 ( .INP(g45), .Z(g4108) );
  INVX0 U1578 ( .INP(n942), .ZN(g4109) );
  INVX0 U1579 ( .INP(g46), .ZN(n942) );
  INVX0 U1580 ( .INP(n940), .ZN(g4112) );
  INVX0 U1581 ( .INP(g47), .ZN(n940) );
  INVX0 U1582 ( .INP(n938), .ZN(g4422) );
  INVX0 U1583 ( .INP(g564), .ZN(n938) );
  NBUFFX2 U1584 ( .INP(g705), .Z(g3222) );
  NBUFFX2 U1585 ( .INP(g43), .Z(g5137) );
  NBUFFX2 U1586 ( .INP(g668), .Z(g5469) );
  NBUFFX2 U1587 ( .INP(g485), .Z(g5468) );
  NOR2X0 U1588 ( .IN1(n69), .IN2(n145), .QN(n550) );
  AO222X1 U1589 ( .IN1(n749), .IN2(n296), .IN3(n297), .IN4(n1026), .IN5(n826), 
        .IN6(g332), .Q(g6795) );
  NAND2X0 U1590 ( .IN1(g277), .IN2(g276), .QN(n333) );
  INVX0 U1591 ( .INP(n235), .ZN(n145) );
  NOR2X0 U1592 ( .IN1(n604), .IN2(g631), .QN(n603) );
  INVX0 U1593 ( .INP(n949), .ZN(n950) );
  INVX0 U1594 ( .INP(n949), .ZN(n951) );
  NAND2X0 U1595 ( .IN1(n178), .IN2(n903), .QN(n656) );
  NOR2X0 U1596 ( .IN1(n893), .IN2(g622), .QN(n629) );
  NAND2X0 U1597 ( .IN1(n832), .IN2(n888), .QN(n192) );
  INVX0 U1598 ( .INP(g102), .ZN(n141) );
  INVX0 U1599 ( .INP(g693), .ZN(n952) );
  INVX0 U1600 ( .INP(g692), .ZN(n954) );
  NOR2X0 U1601 ( .IN1(n674), .IN2(g578), .QN(n482) );
  AO22X1 U1602 ( .IN1(n1041), .IN2(n953), .IN3(n557), .IN4(n992), .Q(g5628) );
  NAND2X0 U1603 ( .IN1(n820), .IN2(n523), .QN(n521) );
  NOR2X0 U1604 ( .IN1(n74), .IN2(n326), .QN(n312) );
  OA21X1 U1605 ( .IN1(n789), .IN2(g207), .IN3(n849), .Q(n565) );
  NOR2X0 U1606 ( .IN1(n59), .IN2(n568), .QN(n556) );
  NOR2X0 U1607 ( .IN1(n624), .IN2(g625), .QN(n623) );
  INVX0 U1608 ( .INP(n957), .ZN(n956) );
  INVX0 U1609 ( .INP(n379), .ZN(n957) );
  NOR2X0 U1610 ( .IN1(g628), .IN2(n613), .QN(n612) );
  NOR2X0 U1611 ( .IN1(n113), .IN2(n561), .QN(n553) );
  INVX0 U1612 ( .INP(n837), .ZN(n959) );
  NOR2X0 U1613 ( .IN1(n339), .IN2(n82), .QN(n323) );
  NOR2X0 U1614 ( .IN1(n322), .IN2(n480), .QN(n339) );
  NOR2X0 U1615 ( .IN1(g582), .IN2(n477), .QN(n476) );
  OA221X1 U1616 ( .IN1(g465), .IN2(n480), .IN3(n481), .IN4(n27), .IN5(n960), 
        .Q(n479) );
  NOR2X0 U1617 ( .IN1(g619), .IN2(n647), .QN(n646) );
  NAND2X0 U1618 ( .IN1(n898), .IN2(n1035), .QN(n283) );
  NAND2X0 U1619 ( .IN1(g697), .IN2(n214), .QN(n209) );
  INVX0 U1620 ( .INP(n864), .ZN(n963) );
  NOR2X0 U1621 ( .IN1(n869), .IN2(n699), .QN(n406) );
  NOR2X0 U1622 ( .IN1(n88), .IN2(n468), .QN(n469) );
  NAND2X0 U1623 ( .IN1(g586), .IN2(n473), .QN(n468) );
  INVX0 U1624 ( .INP(g598), .ZN(n964) );
  INVX0 U1625 ( .INP(n879), .ZN(n967) );
  INVX0 U1626 ( .INP(n963), .ZN(n6) );
  INVX0 U1627 ( .INP(n839), .ZN(n969) );
  INVX0 U1628 ( .INP(n839), .ZN(n970) );
  INVX0 U1629 ( .INP(n715), .ZN(n971) );
  INVX0 U1630 ( .INP(n838), .ZN(n973) );
  NAND2X0 U1631 ( .IN1(n167), .IN2(n921), .QN(n628) );
  NAND2X0 U1632 ( .IN1(n794), .IN2(n921), .QN(n190) );
  NAND2X0 U1633 ( .IN1(n697), .IN2(n921), .QN(n186) );
  OA21X1 U1634 ( .IN1(n922), .IN2(g594), .IN3(n29), .Q(g6304) );
  NAND2X0 U1635 ( .IN1(n895), .IN2(n465), .QN(g6437) );
  NAND2X0 U1636 ( .IN1(n895), .IN2(n467), .QN(g6426) );
  INVX0 U1637 ( .INP(n474), .ZN(n29) );
  NAND2X0 U1638 ( .IN1(n508), .IN2(n758), .QN(n506) );
  NAND2X0 U1639 ( .IN1(g135), .IN2(n618), .QN(n620) );
  NOR2X0 U1640 ( .IN1(g128), .IN2(g131), .QN(n618) );
  NOR2X0 U1641 ( .IN1(n651), .IN2(g616), .QN(n652) );
  INVX0 U1642 ( .INP(g684), .ZN(n57) );
  AO22X1 U1643 ( .IN1(n1036), .IN2(n755), .IN3(n989), .IN4(n279), .Q(n276) );
  INVX0 U1644 ( .INP(n847), .ZN(n977) );
  INVX0 U1645 ( .INP(g690), .ZN(n980) );
  INVX0 U1646 ( .INP(n980), .ZN(n981) );
  NOR2X0 U1647 ( .IN1(n105), .IN2(n650), .QN(n651) );
  NAND2X0 U1648 ( .IN1(n128), .IN2(n487), .QN(n471) );
  NAND2X0 U1649 ( .IN1(n138), .IN2(n819), .QN(n547) );
  NAND2X0 U1650 ( .IN1(g114), .IN2(n618), .QN(n621) );
  NOR2X0 U1651 ( .IN1(g602), .IN2(n870), .QN(g2861) );
  NAND2X0 U1652 ( .IN1(g610), .IN2(g602), .QN(n650) );
  INVX0 U1653 ( .INP(n1038), .ZN(n982) );
  NOR2X0 U1654 ( .IN1(n232), .IN2(n171), .QN(n176) );
  INVX0 U1655 ( .INP(g567), .ZN(n984) );
  INVX0 U1656 ( .INP(n984), .ZN(n985) );
  INVX0 U1657 ( .INP(n171), .ZN(n85) );
  NAND2X0 U1658 ( .IN1(n867), .IN2(n549), .QN(n540) );
  INVX0 U1659 ( .INP(g197), .ZN(n988) );
  INVX0 U1660 ( .INP(n988), .ZN(n989) );
  INVX0 U1661 ( .INP(n988), .ZN(n990) );
  INVX0 U1662 ( .INP(n1040), .ZN(n992) );
  AO221X1 U1663 ( .IN1(n249), .IN2(n250), .IN3(n251), .IN4(n252), .IN5(n1010), 
        .Q(n248) );
  NAND2X0 U1664 ( .IN1(n1045), .IN2(n79), .QN(g6176) );
  NAND2X0 U1665 ( .IN1(n1046), .IN2(n127), .QN(g6179) );
  NAND2X0 U1666 ( .IN1(n1044), .IN2(n118), .QN(g6182) );
  NAND2X0 U1667 ( .IN1(g301), .IN2(n790), .QN(n239) );
  NAND2X0 U1668 ( .IN1(n300), .IN2(n790), .QN(n625) );
  NAND2X0 U1669 ( .IN1(n805), .IN2(n790), .QN(n242) );
  NOR2X0 U1670 ( .IN1(n995), .IN2(n1030), .QN(n994) );
  AO22X1 U1671 ( .IN1(g5627), .IN2(n979), .IN3(g5624), .IN4(n876), .Q(n995) );
  NAND2X0 U1672 ( .IN1(n1044), .IN2(n50), .QN(g6173) );
  OAI221X1 U1673 ( .IN1(n271), .IN2(n112), .IN3(n41), .IN4(n272), .IN5(n990), 
        .QN(n1001) );
  NBUFFX2 U1674 ( .INP(n87), .Z(n1040) );
  NOR3X0 U1675 ( .IN1(n997), .IN2(n998), .IN3(n999), .QN(n996) );
  AO22X1 U1676 ( .IN1(g5628), .IN2(n978), .IN3(g5626), .IN4(n876), .Q(n997) );
  AO222X1 U1677 ( .IN1(n865), .IN2(g414), .IN3(n24), .IN4(g512), .IN5(n855), 
        .IN6(g449), .Q(n999) );
  NAND4X0 U1678 ( .IN1(n1002), .IN2(n1001), .IN3(n1003), .IN4(n1004), .QN(
        n1007) );
  AND2X1 U1679 ( .IN1(n273), .IN2(n274), .Q(n1002) );
  OAI221X1 U1680 ( .IN1(n63), .IN2(n271), .IN3(n710), .IN4(n272), .IN5(n1017), 
        .QN(n1003) );
  OAI222X1 U1681 ( .IN1(n990), .IN2(n110), .IN3(g337), .IN4(n260), .IN5(n266), 
        .IN6(n1036), .QN(n1004) );
  AO22X1 U1682 ( .IN1(n1007), .IN2(n1006), .IN3(n1008), .IN4(n1005), .Q(n1020)
         );
  OAI221X1 U1683 ( .IN1(n260), .IN2(n1040), .IN3(n94), .IN4(n261), .IN5(n977), 
        .QN(n1008) );
  NBUFFX2 U1684 ( .INP(n1017), .Z(n1009) );
  NBUFFX2 U1685 ( .INP(n993), .Z(n1010) );
  NBUFFX2 U1686 ( .INP(n1039), .Z(n1011) );
  NAND2X0 U1687 ( .IN1(g49), .IN2(n447), .QN(n446) );
  INVX0 U1688 ( .INP(g323), .ZN(n71) );
  INVX0 U1689 ( .INP(n120), .ZN(n1037) );
  NOR2X0 U1690 ( .IN1(g310), .IN2(g306), .QN(n455) );
  NAND2X0 U1691 ( .IN1(n1046), .IN2(n84), .QN(g6189) );
  INVX0 U1692 ( .INP(g6794), .ZN(n1018) );
  INVX0 U1693 ( .INP(n1018), .ZN(n1019) );
  NBUFFX2 U1694 ( .INP(n123), .Z(n1036) );
  AND2X1 U1695 ( .IN1(n1020), .IN2(n1021), .Q(n247) );
  AO221X1 U1696 ( .IN1(n251), .IN2(g681), .IN3(n249), .IN4(g679), .IN5(n992), 
        .Q(n1021) );
  INVX0 U1697 ( .INP(n791), .ZN(n1022) );
  INVX0 U1698 ( .INP(n155), .ZN(n1027) );
  INVX0 U1699 ( .INP(g41), .ZN(n155) );
  INVX0 U1700 ( .INP(n989), .ZN(n123) );
  OA21X1 U1701 ( .IN1(n560), .IN2(g279), .IN3(n561), .Q(n558) );
  NOR2X0 U1702 ( .IN1(n87), .IN2(n552), .QN(n551) );
  INVX0 U1703 ( .INP(g269), .ZN(n87) );
  AOI221X1 U1704 ( .IN1(n406), .IN2(n1012), .IN3(n407), .IN4(n56), .IN5(n896), 
        .QN(n1028) );
  NAND2X1 U1705 ( .IN1(n368), .IN2(n994), .QN(g6481) );
  NAND2X1 U1706 ( .IN1(n996), .IN2(n361), .QN(g6482) );
  NOR2X0 U1707 ( .IN1(n862), .IN2(n156), .QN(g3814) );
  NAND2X1 U1708 ( .IN1(n366), .IN2(n367), .QN(n1030) );
  INVX0 U1709 ( .INP(n284), .ZN(n3) );
  NAND2X0 U1710 ( .IN1(n685), .IN2(n434), .QN(n433) );
  NOR2X0 U1711 ( .IN1(n704), .IN2(n592), .QN(n590) );
  NAND2X0 U1712 ( .IN1(g378), .IN2(n407), .QN(n435) );
  NAND2X0 U1713 ( .IN1(g374), .IN2(n407), .QN(n442) );
  INVX0 U1714 ( .INP(n763), .ZN(n1043) );
  NAND2X0 U1715 ( .IN1(g345), .IN2(n593), .QN(n595) );
  NAND2X0 U1716 ( .IN1(g323), .IN2(n593), .QN(n596) );
  NOR2X0 U1717 ( .IN1(n145), .IN2(n1026), .QN(n299) );
  NOR2X0 U1718 ( .IN1(n431), .IN2(n894), .QN(n430) );
  NOR2X0 U1719 ( .IN1(n419), .IN2(n894), .QN(n418) );
  NOR2X0 U1720 ( .IN1(n426), .IN2(n896), .QN(n425) );
  NOR2X0 U1721 ( .IN1(n711), .IN2(n85), .QN(n260) );
  INVX0 U1722 ( .INP(n394), .ZN(n86) );
endmodule

