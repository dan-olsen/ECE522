
module dff_test_0 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_1 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_2 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_3 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_4 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_5 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_6 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_7 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_8 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_9 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_10 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_11 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_12 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_13 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module s298 ( CK, G0, G1, G117, G118, G132, G133, G2, G66, G67, test_si, 
        test_so, test_se );
  input CK, G0, G1, G2, test_si, test_se;
  output G117, G118, G132, G133, G66, G67, test_so;
  wire   G10, G29, G11, G30, G12, G34, G13, G39, G14, G44, G15, G56, G16, G86,
         G17, G92, G18, G98, G19, G102, G20, G107, G21, G113, G22, G119, G23,
         G125, n84, n85, n86, n87, n88, n89, n90, n91, n93, n94, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n185, n186, n187, n188, n189;
  assign G66 = G16;
  assign G67 = G17;
  assign G117 = G18;
  assign G118 = G19;
  assign G132 = G20;
  assign G133 = G21;

  dff_test_13 DFF_0 ( .CK(CK), .Q(G10), .D(G29), .test_si(test_si), .test_so(
        n183), .test_se(n186) );
  dff_test_0 DFF_1 ( .CK(CK), .Q(G11), .D(G30), .test_si(n183), .test_so(n182), 
        .test_se(n187) );
  dff_test_1 DFF_2 ( .CK(CK), .Q(G12), .D(G34), .test_si(n182), .test_so(n181), 
        .test_se(n188) );
  dff_test_2 DFF_3 ( .CK(CK), .Q(G13), .D(G39), .test_si(n181), .test_so(n180), 
        .test_se(n189) );
  dff_test_3 DFF_4 ( .CK(CK), .Q(G14), .D(G44), .test_si(n180), .test_so(n179), 
        .test_se(n186) );
  dff_test_4 DFF_5 ( .CK(CK), .Q(G15), .D(G56), .test_si(n179), .test_so(n178), 
        .test_se(n187) );
  dff_test_5 DFF_6 ( .CK(CK), .Q(G16), .D(G86), .test_si(n178), .test_so(n177), 
        .test_se(n188) );
  dff_test_6 DFF_7 ( .CK(CK), .Q(G17), .D(G92), .test_si(n177), .test_so(n176), 
        .test_se(n189) );
  dff_test_7 DFF_8 ( .CK(CK), .Q(G18), .D(G98), .test_si(n176), .test_so(n175), 
        .test_se(n186) );
  dff_test_8 DFF_9 ( .CK(CK), .Q(G19), .D(G102), .test_si(n175), .test_so(n174), .test_se(n187) );
  dff_test_9 DFF_10 ( .CK(CK), .Q(G20), .D(G107), .test_si(n174), .test_so(
        n173), .test_se(n188) );
  dff_test_10 DFF_11 ( .CK(CK), .Q(G21), .D(G113), .test_si(n173), .test_so(
        n172), .test_se(n189) );
  dff_test_11 DFF_12 ( .CK(CK), .Q(G22), .D(G119), .test_si(n172), .test_so(
        n171), .test_se(n186) );
  dff_test_12 DFF_13 ( .CK(CK), .Q(G23), .D(G125), .test_si(n171), .test_so(
        test_so), .test_se(n187) );
  NOR4X1 U74 ( .IN1(n163), .IN2(n165), .IN3(n119), .IN4(n120), .QN(G34) );
  AO21X1 U106 ( .IN1(n103), .IN2(n157), .IN3(G18), .Q(n100) );
  OAI222X1 U108 ( .IN1(n137), .IN2(n166), .IN3(n91), .IN4(n107), .IN5(n103), 
        .IN6(n137), .QN(n104) );
  OA221X1 U109 ( .IN1(n152), .IN2(n146), .IN3(G16), .IN4(n142), .IN5(n108), 
        .Q(G86) );
  AND4X1 U110 ( .IN1(n99), .IN2(n113), .IN3(n114), .IN4(n112), .Q(G44) );
  NAND4X0 U111 ( .IN1(n151), .IN2(n168), .IN3(n165), .IN4(n152), .QN(n113) );
  XNOR2X1 U114 ( .IN1(n167), .IN2(n119), .Q(n118) );
  XNOR2X1 U118 ( .IN1(G23), .IN2(G1), .Q(n124) );
  XNOR2X1 U119 ( .IN1(G22), .IN2(G2), .Q(n125) );
  AOI22X1 U120 ( .IN1(n143), .IN2(n142), .IN3(G21), .IN4(n146), .QN(n126) );
  OA221X1 U121 ( .IN1(n106), .IN2(G20), .IN3(n141), .IN4(n144), .IN5(n168), 
        .Q(n127) );
  AND3X1 U122 ( .IN1(n129), .IN2(n128), .IN3(n130), .Q(G102) );
  OA22X1 U125 ( .IN1(n103), .IN2(n97), .IN3(n90), .IN4(n142), .Q(n131) );
  INVX0 U128 ( .INP(n155), .ZN(n143) );
  NAND3X0 U129 ( .IN1(n142), .IN2(n98), .IN3(n116), .QN(n112) );
  NBUFFX2 U130 ( .INP(n115), .Z(n161) );
  OR3X1 U131 ( .IN1(G22), .IN2(n155), .IN3(G12), .Q(n138) );
  INVX0 U132 ( .INP(n156), .ZN(n141) );
  NAND3X1 U133 ( .IN1(n102), .IN2(n157), .IN3(n131), .QN(n129) );
  OR2X1 U134 ( .IN1(n132), .IN2(n153), .Q(n134) );
  AO21X1 U135 ( .IN1(n167), .IN2(n91), .IN3(n164), .Q(n123) );
  INVX0 U136 ( .INP(n144), .ZN(n132) );
  NAND3X0 U137 ( .IN1(n132), .IN2(n155), .IN3(n146), .QN(n101) );
  AND3X1 U138 ( .IN1(n146), .IN2(n152), .IN3(n97), .Q(n133) );
  AND2X1 U139 ( .IN1(n135), .IN2(n84), .Q(G29) );
  DELLN1X2 U140 ( .INP(G10), .Z(n151) );
  INVX0 U141 ( .INP(G0), .ZN(n135) );
  INVX0 U142 ( .INP(n135), .ZN(n136) );
  NAND3X1 U143 ( .IN1(n161), .IN2(n167), .IN3(G10), .QN(n116) );
  INVX0 U144 ( .INP(G13), .ZN(n166) );
  NBUFFX2 U145 ( .INP(G17), .Z(n137) );
  NAND3X0 U146 ( .IN1(n105), .IN2(n115), .IN3(G22), .QN(n110) );
  INVX0 U147 ( .INP(n153), .ZN(n139) );
  INVX0 U148 ( .INP(n93), .ZN(n153) );
  INVX0 U149 ( .INP(G14), .ZN(n145) );
  NOR3X0 U150 ( .IN1(n150), .IN2(n126), .IN3(n134), .QN(G113) );
  NAND2X0 U151 ( .IN1(n149), .IN2(n133), .QN(n130) );
  INVX0 U152 ( .INP(n91), .ZN(n140) );
  NOR2X0 U153 ( .IN1(n156), .IN2(G12), .QN(n115) );
  INVX0 U154 ( .INP(G11), .ZN(n155) );
  NOR2X0 U155 ( .IN1(n93), .IN2(n138), .QN(n111) );
  INVX0 U156 ( .INP(n159), .ZN(n91) );
  INVX0 U157 ( .INP(G29), .ZN(n85) );
  OA22X1 U158 ( .IN1(n141), .IN2(n85), .IN3(n84), .IN4(n123), .Q(n122) );
  NBUFFX2 U159 ( .INP(G14), .Z(n147) );
  INVX0 U160 ( .INP(n162), .ZN(n163) );
  INVX0 U161 ( .INP(n110), .ZN(n89) );
  INVX0 U162 ( .INP(n101), .ZN(n87) );
  NAND2X1 U163 ( .IN1(G23), .IN2(n146), .QN(n114) );
  NOR2X0 U164 ( .IN1(n163), .IN2(n124), .QN(G125) );
  INVX0 U165 ( .INP(G23), .ZN(n98) );
  INVX0 U166 ( .INP(G19), .ZN(n97) );
  INVX0 U167 ( .INP(n158), .ZN(n159) );
  INVX0 U168 ( .INP(n144), .ZN(n106) );
  INVX0 U169 ( .INP(G12), .ZN(n158) );
  NOR2X0 U170 ( .IN1(n163), .IN2(n125), .QN(G119) );
  OA21X1 U171 ( .IN1(n136), .IN2(n165), .IN3(n85), .Q(n117) );
  INVX0 U172 ( .INP(n164), .ZN(n99) );
  OAI21X1 U173 ( .IN1(G15), .IN2(n89), .IN3(n148), .QN(n154) );
  NBUFFX2 U174 ( .INP(n86), .Z(n160) );
  OR2X1 U175 ( .IN1(n154), .IN2(n84), .Q(n128) );
  NBUFFX2 U176 ( .INP(n145), .Z(n142) );
  AND2X1 U177 ( .IN1(n148), .IN2(G15), .Q(n109) );
  INVX0 U178 ( .INP(G15), .ZN(n96) );
  NOR4X0 U179 ( .IN1(n150), .IN2(n87), .IN3(n104), .IN4(n153), .QN(G92) );
  AO21X1 U180 ( .IN1(n96), .IN2(n110), .IN3(n111), .Q(n102) );
  NAND2X0 U181 ( .IN1(n158), .IN2(n94), .QN(n144) );
  INVX0 U182 ( .INP(n86), .ZN(n149) );
  INVX0 U183 ( .INP(n145), .ZN(n146) );
  INVX0 U184 ( .INP(n111), .ZN(n148) );
  INVX0 U185 ( .INP(n154), .ZN(n150) );
  NBUFFX2 U186 ( .INP(n147), .Z(n168) );
  AND4X1 U187 ( .IN1(n100), .IN2(n101), .IN3(n149), .IN4(n139), .Q(G98) );
  INVX0 U188 ( .INP(n166), .ZN(n152) );
  INVX0 U189 ( .INP(n166), .ZN(n167) );
  NOR2X0 U190 ( .IN1(n121), .IN2(n122), .QN(G30) );
  AND2X1 U191 ( .IN1(n121), .IN2(n159), .Q(n119) );
  NOR2X0 U192 ( .IN1(n94), .IN2(n147), .QN(n105) );
  NOR2X0 U193 ( .IN1(n117), .IN2(n118), .QN(G39) );
  INVX0 U194 ( .INP(n88), .ZN(n156) );
  INVX0 U195 ( .INP(n152), .ZN(n157) );
  INVX0 U196 ( .INP(n105), .ZN(n93) );
  NOR2X0 U197 ( .IN1(n84), .IN2(n141), .QN(n121) );
  INVX0 U198 ( .INP(G13), .ZN(n94) );
  OA21X1 U199 ( .IN1(n109), .IN2(n89), .IN3(n99), .Q(G56) );
  INVX0 U200 ( .INP(n102), .ZN(n86) );
  INVX0 U201 ( .INP(G10), .ZN(n84) );
  INVX0 U202 ( .INP(G11), .ZN(n88) );
  NAND2X0 U203 ( .IN1(n143), .IN2(n142), .QN(n107) );
  INVX0 U204 ( .INP(G0), .ZN(n162) );
  INVX0 U205 ( .INP(n162), .ZN(n164) );
  INVX0 U206 ( .INP(n90), .ZN(n165) );
  INVX0 U207 ( .INP(n161), .ZN(n90) );
  OA21X1 U208 ( .IN1(n160), .IN2(n127), .IN3(n128), .Q(G107) );
  NOR2X0 U209 ( .IN1(n160), .IN2(n132), .QN(n108) );
  NOR2X0 U210 ( .IN1(n151), .IN2(n140), .QN(n120) );
  NAND2X0 U211 ( .IN1(n159), .IN2(n168), .QN(n103) );
  IBUFFX16 U212 ( .INP(test_se), .ZN(n185) );
  IBUFFX16 U213 ( .INP(n185), .ZN(n186) );
  IBUFFX16 U214 ( .INP(n185), .ZN(n187) );
  IBUFFX16 U215 ( .INP(n185), .ZN(n188) );
  IBUFFX16 U216 ( .INP(n185), .ZN(n189) );
endmodule

