
module dff_test_0 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_1 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_2 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_3 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_4 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_5 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n2;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n2) );
  INVX0 U3 ( .INP(n2), .ZN(Q) );
endmodule


module dff_test_6 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_7 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_8 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n2;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n2) );
  INVX0 U3 ( .INP(n2), .ZN(Q) );
endmodule


module dff_test_9 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_10 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_11 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_12 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_13 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_14 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_15 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_16 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_17 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_18 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_19 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_20 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_21 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_22 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_23 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_24 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_25 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_26 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_27 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_28 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_29 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_30 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_31 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_32 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_33 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_34 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_35 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_36 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_37 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_38 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_39 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_40 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_41 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_42 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n3;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n3) );
  INVX0 U3 ( .INP(n3), .ZN(Q) );
endmodule


module dff_test_43 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_44 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_45 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_46 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_47 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_48 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_49 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_50 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_51 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_52 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_53 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_54 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_55 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_56 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_57 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_58 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_59 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_60 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_61 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_62 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_63 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_64 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_65 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_66 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_67 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_68 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_69 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_70 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_71 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_72 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_73 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_74 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_75 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_76 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_77 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_78 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_79 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_80 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_81 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_82 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_83 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_84 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_85 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_86 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_87 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_88 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_89 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_90 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_91 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n2;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n2) );
  INVX0 U3 ( .INP(n2), .ZN(Q) );
endmodule


module dff_test_92 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_93 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_94 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_95 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_96 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_97 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n3;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n3) );
  INVX0 U3 ( .INP(n3), .ZN(Q) );
endmodule


module dff_test_98 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_99 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_100 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_101 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_102 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_103 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_104 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_105 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_106 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n2;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n2) );
  INVX1 U3 ( .INP(n2), .ZN(Q) );
endmodule


module dff_test_107 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_108 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_109 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_110 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_111 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_112 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_113 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_114 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_115 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_116 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n2;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n2) );
  INVX0 U3 ( .INP(n2), .ZN(Q) );
endmodule


module dff_test_117 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_118 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_119 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_120 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_121 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_122 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n3;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n3) );
  INVX1 U3 ( .INP(n3), .ZN(Q) );
endmodule


module dff_test_123 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_124 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_125 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_126 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_127 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n2;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n2) );
  INVX0 U3 ( .INP(n2), .ZN(Q) );
endmodule


module dff_test_128 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_129 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_130 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_131 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_132 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_133 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_134 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_135 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_136 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_137 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_138 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_139 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_140 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_141 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_142 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_143 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_144 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_145 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_146 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_147 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_148 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_149 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_150 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_151 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_152 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_153 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_154 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_155 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_156 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_157 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_158 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_159 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_160 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_161 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_162 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_163 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_164 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_165 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_166 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_167 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_168 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n2;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n2) );
  INVX0 U3 ( .INP(n2), .ZN(Q) );
endmodule


module dff_test_169 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_170 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_171 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_172 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_173 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_174 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_175 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_176 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_177 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n2;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n2) );
  INVX0 U3 ( .INP(n2), .ZN(Q) );
endmodule


module dff_test_178 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_179 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_180 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_181 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_182 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_183 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_184 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_185 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_186 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_187 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_188 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_189 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_190 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n2;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n2) );
  INVX0 U3 ( .INP(n2), .ZN(Q) );
endmodule


module dff_test_191 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_192 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_193 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_194 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_195 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_196 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_197 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_198 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_199 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_200 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;
  wire   n2;

  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(test_so), 
        .QN(n2) );
  INVX0 U3 ( .INP(n2), .ZN(Q) );
endmodule


module dff_test_201 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_202 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_203 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_204 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_205 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_206 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_207 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_208 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_209 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module dff_test_210 ( CK, Q, D, test_si, test_so, test_se );
  input CK, D, test_si, test_se;
  output Q, test_so;


  SDFFX1 Q_reg ( .D(D), .SI(test_si), .SE(test_se), .CLK(CK), .Q(Q), .QN(
        test_so) );
endmodule


module s9234 ( CK, g102, g107, g1290, g1293, g22, g23, g2584, g301, g306, g310, 
        g314, g319, g32, g3222, g36, g3600, g37, g38, g39, g40, g4098, g4099, 
        g41, g4100, g4101, g4102, g4103, g4104, g4105, g4106, g4107, g4108, 
        g4109, g4110, g4112, g4121, g42, g4307, g4321, g44, g4422, g45, g46, 
        g47, g4809, g5137, g5468, g5469, g557, g558, g559, g560, g561, g562, 
        g563, g564, g567, g5692, g6282, g6284, g6360, g6362, g6364, g6366, 
        g6368, g6370, g6372, g6374, g639, g6728, g702, g705, g89, g94, g98, 
        test_si, test_so, test_se );
  input CK, g102, g107, g22, g23, g301, g306, g310, g314, g319, g32, g36, g37,
         g38, g39, g40, g41, g42, g44, g45, g46, g47, g557, g558, g559, g560,
         g561, g562, g563, g564, g567, g639, g702, g705, g89, g94, g98,
         test_si, test_se;
  output g1290, g1293, g2584, g3222, g3600, g4098, g4099, g4100, g4101, g4102,
         g4103, g4104, g4105, g4106, g4107, g4108, g4109, g4110, g4112, g4121,
         g4307, g4321, g4422, g4809, g5137, g5468, g5469, g5692, g6282, g6284,
         g6360, g6362, g6364, g6366, g6368, g6370, g6372, g6374, g6728,
         test_so;
  wire   g678, g332, g123, g207, g695, g461, g18, g292, g331, g689, g24, g465,
         g84, g291, g676, g622, g117, g278, g128, g598, g554, g496, g179, g48,
         g590, g551, g682, g606, g188, g646, g327, g361, g289, g398, g5700,
         g684, g619, g208, g248, g390, g5698, g625, g681, g437, g276, g323,
         g224, g685, g157, g5470, g282, g697, g206, g449, g118, g528, g284,
         g426, g634, g669, g520, g281, g175, g5472, g631, g69, g693, g337,
         g457, g486, g471, g328, g285, g418, g402, g297, g212, g410, g430,
         g662, g453, g269, g574, g441, g664, g349, g211, g586, g571, g326,
         g698, g654, g293, g690, g445, g374, g5694, g6, g687, g357, g386,
         g5697, g504, g665, g166, g5471, g541, g74, g338, g696, g516, g536,
         g683, g353, g545, g254, g341, g290, g2, g287, g336, g345, g628, g679,
         g28, g688, g283, g613, g10, g14, g680, g143, g672, g667, g366, g279,
         g492, g170, g686, g288, g638, g602, g642, g280, g663, g610, g148,
         g209, g675, g478, g122, g54, g594, g286, g489, g616, g79, g218, g242,
         g578, g184, g5473, g119, g139, g422, g210, g394, g5699, g230, g204,
         g658, g650, g378, g5695, g508, g548, g370, g5693, g406, g236, g500,
         g205, g197, g666, g114, g524, g260, g111, g131, g677, g582, g193,
         g5474, g135, g382, g5696, g414, g434, g266, g49, g152, g692, g277,
         g127, g161, g512, g532, g64, g694, g691, g1, g59, g5624, g6294, g5386,
         g6688, g6110, g6300, g6485, g4757, g6173, g6182, g6426, g4430, g2859,
         g6795, g6686, g3725, g4446, g6292, g6689, g6481, g6297, g5231, g5531,
         g3729, g5626, g4447, g3731, g2670, g6293, g6690, g6179, g6791, g6691,
         g6794, g6453, g6113, g6167, g4444, g5627, g6792, g6286, g6684, g4740,
         g6109, g4458, g6307, g4454, g5916, g5628, g3727, g6455, g5291, g4433,
         g6845, g6483, g4219, g6176, g3724, g6299, g6142, g6704, g4752, g6309,
         g6787, g6454, g6456, g4872, g4497, g6296, g5625, g4460, g3768, g6793,
         g4607, g4501, g4440, g6790, g6452, g6185, g4436, g3828, g6310, g6687,
         g5629, g6937, g3454, g6921, g6301, g5532, g4441, g4157, g3730, g5303,
         g5533, g6170, g5277, g4443, g6304, g6844, g6189, g6116, g5583, g4761,
         g5535, g5622, g6480, g6447, g6298, g2433, g6290, g6114, g4451, g6685,
         g6450, g6437, g6789, g6291, g5323, g3728, g6444, g5295, g6118, g2861,
         g5050, g4434, g4687, g6108, g6287, g3844, g4438, g1802, g3726, g6482,
         g5017, g3910, g6303, g6440, g5149, g5701, g6788, g6702, g4773, g6936,
         g4450, g3814, g6295, g5167, g4455, g3599, g6289, g6479, n655, n656,
         n2116, n1048, n1050, n1051, n1054, n1055, n1056, n1057, n1058, n1059,
         n1062, n1063, n1064, n1065, n1066, n1069, n1070, n1072, n1073, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1133, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1184, n1185, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1202, n1203, n1204, n1205,
         n1206, n1207, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1493, n1494, n1496, n1497,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1722, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1759, n1760, n1761, n1762,
         n1763, n1765, n1766, n1767, n1768, n1770, n1772, n1774, n1776, n1778,
         n1780, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2339, n2340, n2341, n2342;
  assign g1290 = g666;
  assign g6284 = g6110;
  assign g6370 = g6173;
  assign g6360 = g6182;
  assign g6374 = g6179;
  assign g6364 = g6167;
  assign g6372 = g6176;
  assign g6362 = g6185;
  assign g6368 = g6170;
  assign g6366 = g6189;
  assign g4809 = g2433;
  assign g2584 = g1802;
  assign g4121 = g3599;

  dff_test_210 DFF_0 ( .CK(CK), .Q(g678), .D(n1915), .test_si(test_si), 
        .test_so(n2337), .test_se(n2340) );
  dff_test_0 DFF_1 ( .CK(CK), .Q(g332), .D(g6795), .test_si(n2337), .test_so(
        n2336), .test_se(n2341) );
  dff_test_1 DFF_2 ( .CK(CK), .Q(g123), .D(g6937), .test_si(n2336), .test_so(
        n2335), .test_se(n2340) );
  dff_test_2 DFF_3 ( .CK(CK), .Q(g207), .D(g5626), .test_si(n2335), .test_so(
        n2334), .test_se(n2341) );
  dff_test_3 DFF_4 ( .CK(CK), .Q(g695), .D(g18), .test_si(n2334), .test_so(
        n2333), .test_se(n2340) );
  dff_test_4 DFF_5 ( .CK(CK), .Q(g461), .D(g4440), .test_si(n2333), .test_so(
        n2332), .test_se(n2341) );
  dff_test_5 DFF_6 ( .CK(CK), .Q(g18), .D(g6684), .test_si(n2332), .test_so(
        n2331), .test_se(n2340) );
  dff_test_6 DFF_7 ( .CK(CK), .Q(g292), .D(g571), .test_si(n2331), .test_so(
        n2330), .test_se(n2341) );
  dff_test_7 DFF_8 ( .CK(CK), .Q(g331), .D(g3730), .test_si(n2330), .test_so(
        n2329), .test_se(n2340) );
  dff_test_8 DFF_9 ( .CK(CK), .Q(g689), .D(g4103), .test_si(n2329), .test_so(
        n2328), .test_se(n2341) );
  dff_test_9 DFF_10 ( .CK(CK), .Q(g24), .D(g6685), .test_si(n2328), .test_so(
        n2327), .test_se(n2340) );
  dff_test_10 DFF_11 ( .CK(CK), .Q(g465), .D(g6297), .test_si(n2327), 
        .test_so(n2326), .test_se(n2341) );
  dff_test_11 DFF_12 ( .CK(CK), .Q(g84), .D(g6456), .test_si(n2326), .test_so(
        n2325), .test_se(n2340) );
  dff_test_12 DFF_13 ( .CK(CK), .Q(g291), .D(g654), .test_si(n2325), .test_so(
        n2324), .test_se(n2341) );
  dff_test_13 DFF_14 ( .CK(CK), .Q(g676), .D(n1078), .test_si(n2324), 
        .test_so(n2323), .test_se(n2340) );
  dff_test_14 DFF_15 ( .CK(CK), .Q(g622), .D(g4460), .test_si(n2323), 
        .test_so(n2322), .test_se(n2341) );
  dff_test_15 DFF_16 ( .CK(CK), .Q(g117), .D(g4497), .test_si(n2322), 
        .test_so(n2321), .test_se(n2340) );
  dff_test_16 DFF_17 ( .CK(CK), .Q(g278), .D(g5627), .test_si(n2321), 
        .test_so(n2320), .test_se(n2341) );
  dff_test_17 DFF_18 ( .CK(CK), .Q(g128), .D(g4773), .test_si(n2320), 
        .test_so(n2319), .test_se(n2340) );
  dff_test_18 DFF_19 ( .CK(CK), .Q(g598), .D(g2859), .test_si(n2319), 
        .test_so(n2318), .test_se(n2341) );
  dff_test_19 DFF_20 ( .CK(CK), .Q(g554), .D(g6790), .test_si(n2318), 
        .test_so(n2317), .test_se(n2340) );
  dff_test_20 DFF_21 ( .CK(CK), .Q(g496), .D(g6702), .test_si(n2317), 
        .test_so(n2316), .test_se(n2341) );
  dff_test_21 DFF_22 ( .CK(CK), .Q(g179), .D(g6116), .test_si(n2316), 
        .test_so(n2315), .test_se(n2340) );
  dff_test_22 DFF_23 ( .CK(CK), .Q(g48), .D(n1115), .test_si(n2315), .test_so(
        n2314), .test_se(n2341) );
  dff_test_23 DFF_24 ( .CK(CK), .Q(g590), .D(g6437), .test_si(n2314), 
        .test_so(n2313), .test_se(n2340) );
  dff_test_24 DFF_25 ( .CK(CK), .Q(g551), .D(g6789), .test_si(n2313), 
        .test_so(n2312), .test_se(n2341) );
  dff_test_25 DFF_26 ( .CK(CK), .Q(g682), .D(g18), .test_si(n2312), .test_so(
        n2311), .test_se(n2340) );
  dff_test_26 DFF_27 ( .CK(CK), .Q(g6689), .D(g6481), .test_si(n2311), 
        .test_so(n2310), .test_se(n2341) );
  dff_test_27 DFF_28 ( .CK(CK), .Q(g606), .D(g4219), .test_si(n2310), 
        .test_so(n2309), .test_se(n2340) );
  dff_test_28 DFF_29 ( .CK(CK), .Q(g188), .D(g6118), .test_si(n2309), 
        .test_so(n2308), .test_se(n2341) );
  dff_test_29 DFF_30 ( .CK(CK), .Q(g646), .D(g4501), .test_si(n2308), 
        .test_so(n2307), .test_se(n2340) );
  dff_test_30 DFF_31 ( .CK(CK), .Q(g327), .D(g3728), .test_si(n2307), 
        .test_so(n2306), .test_se(n2341) );
  dff_test_31 DFF_32 ( .CK(CK), .Q(g361), .D(g6440), .test_si(n2306), 
        .test_so(n2305), .test_se(n2340) );
  dff_test_32 DFF_33 ( .CK(CK), .Q(g289), .D(g646), .test_si(n2305), .test_so(
        n2304), .test_se(n2341) );
  dff_test_33 DFF_34 ( .CK(CK), .Q(g398), .D(g5700), .test_si(n2304), 
        .test_so(n2303), .test_se(n2340) );
  dff_test_34 DFF_35 ( .CK(CK), .Q(g684), .D(n1923), .test_si(n2303), 
        .test_so(n2302), .test_se(n2341) );
  dff_test_35 DFF_36 ( .CK(CK), .Q(g619), .D(g4157), .test_si(n2302), 
        .test_so(n2301), .test_se(n2340) );
  dff_test_36 DFF_37 ( .CK(CK), .Q(g208), .D(g5533), .test_si(n2301), 
        .test_so(n2300), .test_se(n2341) );
  dff_test_37 DFF_38 ( .CK(CK), .Q(g248), .D(n1800), .test_si(n2300), 
        .test_so(n2299), .test_se(n2340) );
  dff_test_38 DFF_39 ( .CK(CK), .Q(g390), .D(g5698), .test_si(n2299), 
        .test_so(n2298), .test_se(n2341) );
  dff_test_39 DFF_40 ( .CK(CK), .Q(g625), .D(g4687), .test_si(n2298), 
        .test_so(n2297), .test_se(n2340) );
  dff_test_40 DFF_41 ( .CK(CK), .Q(g681), .D(g14), .test_si(n2297), .test_so(
        n2296), .test_se(n2341) );
  dff_test_41 DFF_42 ( .CK(CK), .Q(g437), .D(g4433), .test_si(n2296), 
        .test_so(n2295), .test_se(n2340) );
  dff_test_42 DFF_43 ( .CK(CK), .Q(g276), .D(g5532), .test_si(n2295), 
        .test_so(n2294), .test_se(n2341) );
  dff_test_43 DFF_44 ( .CK(CK), .Q(g6686), .D(g6479), .test_si(n2294), 
        .test_so(n2293), .test_se(n2340) );
  dff_test_44 DFF_45 ( .CK(CK), .Q(g323), .D(g3731), .test_si(n2293), 
        .test_so(n2292), .test_se(n2341) );
  dff_test_45 DFF_46 ( .CK(CK), .Q(g224), .D(n1831), .test_si(n2292), 
        .test_so(n2291), .test_se(n2340) );
  dff_test_46 DFF_47 ( .CK(CK), .Q(g685), .D(g4099), .test_si(n2291), 
        .test_so(n2290), .test_se(n2341) );
  dff_test_47 DFF_48 ( .CK(CK), .Q(g5137), .D(g6142), .test_si(n2290), 
        .test_so(n2289), .test_se(n2340) );
  dff_test_48 DFF_49 ( .CK(CK), .Q(g157), .D(g5470), .test_si(n2289), 
        .test_so(n2288), .test_se(n2341) );
  dff_test_49 DFF_50 ( .CK(CK), .Q(g282), .D(g6793), .test_si(n2288), 
        .test_so(n2287), .test_se(n2340) );
  dff_test_50 DFF_51 ( .CK(CK), .Q(g697), .D(n1923), .test_si(n2287), 
        .test_so(n2286), .test_se(n2341) );
  dff_test_51 DFF_52 ( .CK(CK), .Q(g206), .D(g5624), .test_si(n2286), 
        .test_so(n2285), .test_se(n2340) );
  dff_test_52 DFF_53 ( .CK(CK), .Q(g449), .D(g4450), .test_si(n2285), 
        .test_so(n2284), .test_se(n2341) );
  dff_test_53 DFF_54 ( .CK(CK), .Q(g118), .D(g3724), .test_si(n2284), 
        .test_so(n2283), .test_se(n2340) );
  dff_test_54 DFF_55 ( .CK(CK), .Q(g528), .D(g6286), .test_si(n2283), 
        .test_so(n2282), .test_se(n2341) );
  dff_test_55 DFF_56 ( .CK(CK), .Q(g284), .D(n2049), .test_si(n2282), 
        .test_so(n2281), .test_se(n2340) );
  dff_test_56 DFF_57 ( .CK(CK), .Q(g426), .D(g4458), .test_si(n2281), 
        .test_so(n2280), .test_se(n2341) );
  dff_test_57 DFF_58 ( .CK(CK), .Q(g634), .D(g3454), .test_si(n2280), 
        .test_so(n2279), .test_se(n2340) );
  dff_test_58 DFF_59 ( .CK(CK), .Q(g669), .D(g5386), .test_si(n2279), 
        .test_so(n2278), .test_se(n2341) );
  dff_test_59 DFF_60 ( .CK(CK), .Q(g520), .D(g6309), .test_si(n2278), 
        .test_so(n2277), .test_se(n2340) );
  dff_test_60 DFF_61 ( .CK(CK), .Q(g281), .D(n1072), .test_si(n2277), 
        .test_so(n2276), .test_se(n2341) );
  dff_test_61 DFF_62 ( .CK(CK), .Q(g175), .D(g5472), .test_si(n2276), 
        .test_so(n2275), .test_se(n2340) );
  dff_test_62 DFF_63 ( .CK(CK), .Q(g6690), .D(g6482), .test_si(n2275), 
        .test_so(n2274), .test_se(n2341) );
  dff_test_63 DFF_64 ( .CK(CK), .Q(g631), .D(g5167), .test_si(n2274), 
        .test_so(n2273), .test_se(n2340) );
  dff_test_64 DFF_65 ( .CK(CK), .Q(g69), .D(g6453), .test_si(n2273), .test_so(
        n2272), .test_se(n2341) );
  dff_test_65 DFF_66 ( .CK(CK), .Q(g693), .D(g10), .test_si(n2272), .test_so(
        n2271), .test_se(n2340) );
  dff_test_66 DFF_67 ( .CK(CK), .Q(g337), .D(n1722), .test_si(n2271), 
        .test_so(n2270), .test_se(n2341) );
  dff_test_67 DFF_68 ( .CK(CK), .Q(g457), .D(g4443), .test_si(n2270), 
        .test_so(n2269), .test_se(n2340) );
  dff_test_68 DFF_69 ( .CK(CK), .Q(g486), .D(n1169), .test_si(n2269), 
        .test_so(n2268), .test_se(n2341) );
  dff_test_69 DFF_70 ( .CK(CK), .Q(g471), .D(g664), .test_si(n2268), .test_so(
        n2267), .test_se(n2340) );
  dff_test_70 DFF_71 ( .CK(CK), .Q(g328), .D(g3729), .test_si(n2267), 
        .test_so(n2266), .test_se(n2341) );
  dff_test_71 DFF_72 ( .CK(CK), .Q(g285), .D(n2043), .test_si(n2266), 
        .test_so(n2265), .test_se(n2340) );
  dff_test_72 DFF_73 ( .CK(CK), .Q(g418), .D(g4451), .test_si(n2265), 
        .test_so(n2264), .test_se(n2341) );
  dff_test_73 DFF_74 ( .CK(CK), .Q(g402), .D(g4438), .test_si(n2264), 
        .test_so(n2263), .test_se(n2340) );
  dff_test_74 DFF_75 ( .CK(CK), .Q(g297), .D(g6298), .test_si(n2263), 
        .test_so(n2262), .test_se(n2341) );
  dff_test_75 DFF_76 ( .CK(CK), .Q(g212), .D(n2049), .test_si(n2262), 
        .test_so(n2261), .test_se(n2340) );
  dff_test_76 DFF_77 ( .CK(CK), .Q(g410), .D(g4444), .test_si(n2261), 
        .test_so(n2260), .test_se(n2341) );
  dff_test_77 DFF_78 ( .CK(CK), .Q(g430), .D(g4434), .test_si(n2260), 
        .test_so(n2259), .test_se(n2340) );
  dff_test_78 DFF_79 ( .CK(CK), .Q(g6687), .D(g6845), .test_si(n2259), 
        .test_so(n2258), .test_se(n2341) );
  dff_test_79 DFF_80 ( .CK(CK), .Q(g662), .D(n1219), .test_si(n2258), 
        .test_so(n2257), .test_se(n2340) );
  dff_test_80 DFF_81 ( .CK(CK), .Q(g453), .D(g4446), .test_si(n2257), 
        .test_so(n2256), .test_se(n2341) );
  dff_test_81 DFF_82 ( .CK(CK), .Q(g269), .D(g6290), .test_si(n2256), 
        .test_so(n2255), .test_se(n2340) );
  dff_test_82 DFF_83 ( .CK(CK), .Q(g574), .D(g6426), .test_si(n2255), 
        .test_so(n2254), .test_se(n2341) );
  dff_test_83 DFF_84 ( .CK(CK), .Q(g441), .D(g4430), .test_si(n2254), 
        .test_so(n2253), .test_se(n2340) );
  dff_test_84 DFF_85 ( .CK(CK), .Q(g664), .D(g663), .test_si(n2253), .test_so(
        n2252), .test_se(n2341) );
  dff_test_85 DFF_86 ( .CK(CK), .Q(g349), .D(g5295), .test_si(n2252), 
        .test_so(n2251), .test_se(n2340) );
  dff_test_86 DFF_87 ( .CK(CK), .Q(g211), .D(g6792), .test_si(n2251), 
        .test_so(n2250), .test_se(n2341) );
  dff_test_87 DFF_88 ( .CK(CK), .Q(g586), .D(g6299), .test_si(n2250), 
        .test_so(n2249), .test_se(n2340) );
  dff_test_88 DFF_89 ( .CK(CK), .Q(g571), .D(g5149), .test_si(n2249), 
        .test_so(n2248), .test_se(n2341) );
  dff_test_89 DFF_90 ( .CK(CK), .Q(g6685), .D(g6844), .test_si(n2248), 
        .test_so(n2247), .test_se(n2340) );
  dff_test_90 DFF_91 ( .CK(CK), .Q(g326), .D(g4607), .test_si(n2247), 
        .test_so(n2246), .test_se(n2341) );
  dff_test_91 DFF_92 ( .CK(CK), .Q(g698), .D(g4105), .test_si(n2246), 
        .test_so(n2245), .test_se(n2340) );
  dff_test_92 DFF_93 ( .CK(CK), .Q(g654), .D(g5017), .test_si(n2245), 
        .test_so(n2244), .test_se(n2341) );
  dff_test_93 DFF_94 ( .CK(CK), .Q(g293), .D(g6294), .test_si(n2244), 
        .test_so(n2243), .test_se(n2340) );
  dff_test_94 DFF_95 ( .CK(CK), .Q(g690), .D(g1), .test_si(n2243), .test_so(
        n2242), .test_se(n2341) );
  dff_test_95 DFF_96 ( .CK(CK), .Q(g445), .D(g4454), .test_si(n2242), 
        .test_so(n2241), .test_se(n2340) );
  dff_test_96 DFF_97 ( .CK(CK), .Q(g374), .D(g5694), .test_si(n2241), 
        .test_so(n2240), .test_se(n2341) );
  dff_test_97 DFF_98 ( .CK(CK), .Q(g6), .D(g6689), .test_si(n2240), .test_so(
        n2239), .test_se(n2340) );
  dff_test_98 DFF_99 ( .CK(CK), .Q(g687), .D(g4101), .test_si(n2239), 
        .test_so(n2238), .test_se(n2341) );
  dff_test_99 DFF_100 ( .CK(CK), .Q(g357), .D(g5303), .test_si(n2238), 
        .test_so(n2237), .test_se(n2340) );
  dff_test_100 DFF_101 ( .CK(CK), .Q(g386), .D(g5697), .test_si(n2237), 
        .test_so(n2236), .test_se(n2341) );
  dff_test_101 DFF_102 ( .CK(CK), .Q(g504), .D(g6296), .test_si(n2236), 
        .test_so(n2235), .test_se(n2340) );
  dff_test_102 DFF_103 ( .CK(CK), .Q(g665), .D(g4106), .test_si(n2235), 
        .test_so(n2234), .test_se(n2341) );
  dff_test_103 DFF_104 ( .CK(CK), .Q(g166), .D(g5471), .test_si(n2234), 
        .test_so(n2233), .test_se(n2340) );
  dff_test_104 DFF_105 ( .CK(CK), .Q(g541), .D(g6289), .test_si(n2233), 
        .test_so(n2232), .test_se(n2341) );
  dff_test_105 DFF_106 ( .CK(CK), .Q(g74), .D(g6454), .test_si(n2232), 
        .test_so(n2231), .test_se(n2340) );
  dff_test_106 DFF_107 ( .CK(CK), .Q(g338), .D(g5323), .test_si(n2231), 
        .test_so(n2230), .test_se(n2341) );
  dff_test_107 DFF_108 ( .CK(CK), .Q(g696), .D(n1912), .test_si(n2230), 
        .test_so(n2229), .test_se(n2340) );
  dff_test_108 DFF_109 ( .CK(CK), .Q(g516), .D(g6307), .test_si(n2229), 
        .test_so(n2228), .test_se(n2341) );
  dff_test_109 DFF_110 ( .CK(CK), .Q(g536), .D(g6293), .test_si(n2228), 
        .test_so(n2227), .test_se(n2340) );
  dff_test_110 DFF_111 ( .CK(CK), .Q(g683), .D(n1912), .test_si(n2227), 
        .test_so(n2226), .test_se(n2341) );
  dff_test_111 DFF_112 ( .CK(CK), .Q(g353), .D(g5050), .test_si(n2226), 
        .test_so(n2225), .test_se(n2340) );
  dff_test_112 DFF_113 ( .CK(CK), .Q(g545), .D(g6787), .test_si(n2225), 
        .test_so(n2224), .test_se(n2341) );
  dff_test_113 DFF_114 ( .CK(CK), .Q(g254), .D(g654), .test_si(n2224), 
        .test_so(n2223), .test_se(n2340) );
  dff_test_114 DFF_115 ( .CK(CK), .Q(g341), .D(g5277), .test_si(n2223), 
        .test_so(n2222), .test_se(n2341) );
  dff_test_115 DFF_116 ( .CK(CK), .Q(g290), .D(n1800), .test_si(n2222), 
        .test_so(n2221), .test_se(n2340) );
  dff_test_116 DFF_117 ( .CK(CK), .Q(g2), .D(g6688), .test_si(n2221), 
        .test_so(n2220), .test_se(n2341) );
  dff_test_117 DFF_118 ( .CK(CK), .Q(g287), .D(g642), .test_si(n2220), 
        .test_so(n2219), .test_se(n2340) );
  dff_test_118 DFF_119 ( .CK(CK), .Q(g336), .D(g6921), .test_si(n2219), 
        .test_so(n2218), .test_se(n2341) );
  dff_test_119 DFF_120 ( .CK(CK), .Q(g345), .D(g5291), .test_si(n2218), 
        .test_so(n2217), .test_se(n2340) );
  dff_test_120 DFF_121 ( .CK(CK), .Q(g628), .D(g4872), .test_si(n2217), 
        .test_so(n2216), .test_se(n2341) );
  dff_test_121 DFF_122 ( .CK(CK), .Q(g679), .D(n1920), .test_si(n2216), 
        .test_so(n2215), .test_se(n2340) );
  dff_test_122 DFF_123 ( .CK(CK), .Q(g28), .D(g6687), .test_si(n2215), 
        .test_so(n2214), .test_se(n2341) );
  dff_test_123 DFF_124 ( .CK(CK), .Q(g688), .D(g4102), .test_si(n2214), 
        .test_so(n2213), .test_se(n2340) );
  dff_test_124 DFF_125 ( .CK(CK), .Q(g283), .D(g6794), .test_si(n2213), 
        .test_so(n2212), .test_se(n2341) );
  dff_test_125 DFF_126 ( .CK(CK), .Q(g613), .D(g3828), .test_si(n2212), 
        .test_so(n2211), .test_se(n2340) );
  dff_test_126 DFF_127 ( .CK(CK), .Q(g10), .D(g6690), .test_si(n2211), 
        .test_so(n2210), .test_se(n2341) );
  dff_test_127 DFF_128 ( .CK(CK), .Q(g14), .D(g6691), .test_si(n2210), 
        .test_so(n2209), .test_se(n2340) );
  dff_test_128 DFF_129 ( .CK(CK), .Q(g680), .D(g10), .test_si(n2209), 
        .test_so(n2208), .test_se(n2341) );
  dff_test_129 DFF_130 ( .CK(CK), .Q(g143), .D(g6108), .test_si(n2208), 
        .test_so(n2207), .test_se(n2340) );
  dff_test_130 DFF_131 ( .CK(CK), .Q(g672), .D(g5231), .test_si(n2207), 
        .test_so(n2206), .test_se(n2341) );
  dff_test_131 DFF_132 ( .CK(CK), .Q(g667), .D(g4108), .test_si(n2206), 
        .test_so(n2205), .test_se(n2340) );
  dff_test_132 DFF_133 ( .CK(CK), .Q(g366), .D(g5916), .test_si(n2205), 
        .test_so(n2204), .test_se(n2341) );
  dff_test_133 DFF_134 ( .CK(CK), .Q(g279), .D(g5628), .test_si(n2204), 
        .test_so(n2203), .test_se(n2340) );
  dff_test_134 DFF_135 ( .CK(CK), .Q(g492), .D(g6704), .test_si(n2203), 
        .test_so(n2202), .test_se(n2341) );
  dff_test_135 DFF_136 ( .CK(CK), .Q(g170), .D(g6114), .test_si(n2202), 
        .test_so(n2201), .test_se(n2340) );
  dff_test_136 DFF_137 ( .CK(CK), .Q(g686), .D(g4100), .test_si(n2201), 
        .test_so(n2200), .test_se(n2341) );
  dff_test_137 DFF_138 ( .CK(CK), .Q(g288), .D(g606), .test_si(n2200), 
        .test_so(n2199), .test_se(n2340) );
  dff_test_138 DFF_139 ( .CK(CK), .Q(g638), .D(g667), .test_si(n2199), 
        .test_so(n2198), .test_se(n2341) );
  dff_test_139 DFF_140 ( .CK(CK), .Q(g602), .D(g2861), .test_si(n2198), 
        .test_so(n2197), .test_se(n2340) );
  dff_test_140 DFF_141 ( .CK(CK), .Q(g642), .D(g3844), .test_si(n2197), 
        .test_so(n2196), .test_se(n2341) );
  dff_test_141 DFF_142 ( .CK(CK), .Q(g280), .D(g5535), .test_si(n2196), 
        .test_so(n2195), .test_se(n2340) );
  dff_test_142 DFF_143 ( .CK(CK), .Q(g663), .D(g4106), .test_si(n2195), 
        .test_so(n2194), .test_se(n2341) );
  dff_test_143 DFF_144 ( .CK(CK), .Q(g610), .D(g2670), .test_si(n2194), 
        .test_so(n2193), .test_se(n2340) );
  dff_test_144 DFF_145 ( .CK(CK), .Q(g148), .D(g5583), .test_si(n2193), 
        .test_so(n2192), .test_se(n2341) );
  dff_test_145 DFF_146 ( .CK(CK), .Q(g209), .D(g5629), .test_si(n2192), 
        .test_so(n2191), .test_se(n2340) );
  dff_test_146 DFF_147 ( .CK(CK), .Q(g675), .D(n1767), .test_si(n2191), 
        .test_so(n2190), .test_se(n2341) );
  dff_test_147 DFF_148 ( .CK(CK), .Q(g478), .D(g665), .test_si(n2190), 
        .test_so(n2189), .test_se(n2340) );
  dff_test_148 DFF_149 ( .CK(CK), .Q(g122), .D(g3726), .test_si(n2189), 
        .test_so(n2188), .test_se(n2341) );
  dff_test_149 DFF_150 ( .CK(CK), .Q(g54), .D(g6447), .test_si(n2188), 
        .test_so(n2187), .test_se(n2340) );
  dff_test_150 DFF_151 ( .CK(CK), .Q(g594), .D(g6304), .test_si(n2187), 
        .test_so(n2186), .test_se(n2341) );
  dff_test_151 DFF_152 ( .CK(CK), .Q(g286), .D(n1830), .test_si(n2186), 
        .test_so(n2185), .test_se(n2340) );
  dff_test_152 DFF_153 ( .CK(CK), .Q(g489), .D(n1987), .test_si(n2185), 
        .test_so(n2184), .test_se(n2341) );
  dff_test_153 DFF_154 ( .CK(CK), .Q(g616), .D(g3768), .test_si(n2184), 
        .test_so(n2183), .test_se(n2340) );
  dff_test_154 DFF_155 ( .CK(CK), .Q(g79), .D(g6455), .test_si(n2183), 
        .test_so(n2182), .test_se(n2341) );
  dff_test_155 DFF_156 ( .CK(CK), .Q(g218), .D(n2043), .test_si(n2182), 
        .test_so(n2181), .test_se(n2340) );
  dff_test_156 DFF_157 ( .CK(CK), .Q(g242), .D(g646), .test_si(n2181), 
        .test_so(n2180), .test_se(n2341) );
  dff_test_157 DFF_158 ( .CK(CK), .Q(g578), .D(g6291), .test_si(n2180), 
        .test_so(n2179), .test_se(n2340) );
  dff_test_158 DFF_159 ( .CK(CK), .Q(g184), .D(g5473), .test_si(n2179), 
        .test_so(n2178), .test_se(n2341) );
  dff_test_159 DFF_160 ( .CK(CK), .Q(g119), .D(g3725), .test_si(n2178), 
        .test_so(n2177), .test_se(n2340) );
  dff_test_160 DFF_161 ( .CK(CK), .Q(g5469), .D(n655), .test_si(n2177), 
        .test_so(n2176), .test_se(n2341) );
  dff_test_161 DFF_162 ( .CK(CK), .Q(g139), .D(g4757), .test_si(n2176), 
        .test_so(n2175), .test_se(n2340) );
  dff_test_162 DFF_163 ( .CK(CK), .Q(g422), .D(g4455), .test_si(n2175), 
        .test_so(n2174), .test_se(n2341) );
  dff_test_163 DFF_164 ( .CK(CK), .Q(g210), .D(g6791), .test_si(n2174), 
        .test_so(n2173), .test_se(n2340) );
  dff_test_164 DFF_165 ( .CK(CK), .Q(g394), .D(g5699), .test_si(n2173), 
        .test_so(n2172), .test_se(n2341) );
  dff_test_165 DFF_166 ( .CK(CK), .Q(g230), .D(g642), .test_si(n2172), 
        .test_so(n2171), .test_se(n2340) );
  dff_test_166 DFF_167 ( .CK(CK), .Q(g6684), .D(g6485), .test_si(n2171), 
        .test_so(n2170), .test_se(n2341) );
  dff_test_167 DFF_168 ( .CK(CK), .Q(g204), .D(g5531), .test_si(n2170), 
        .test_so(n2169), .test_se(n2340) );
  dff_test_168 DFF_169 ( .CK(CK), .Q(g658), .D(g3814), .test_si(n2169), 
        .test_so(n2168), .test_se(n2341) );
  dff_test_169 DFF_170 ( .CK(CK), .Q(g650), .D(g4761), .test_si(n2168), 
        .test_so(n2167), .test_se(n2340) );
  dff_test_170 DFF_171 ( .CK(CK), .Q(g378), .D(g5695), .test_si(n2167), 
        .test_so(n2166), .test_se(n2341) );
  dff_test_171 DFF_172 ( .CK(CK), .Q(g508), .D(g6300), .test_si(n2166), 
        .test_so(n2165), .test_se(n2340) );
  dff_test_172 DFF_173 ( .CK(CK), .Q(g548), .D(g6788), .test_si(n2165), 
        .test_so(n2164), .test_se(n2341) );
  dff_test_173 DFF_174 ( .CK(CK), .Q(g370), .D(g5693), .test_si(n2164), 
        .test_so(n2163), .test_se(n2340) );
  dff_test_174 DFF_175 ( .CK(CK), .Q(g406), .D(g4441), .test_si(n2163), 
        .test_so(n2162), .test_se(n2341) );
  dff_test_175 DFF_176 ( .CK(CK), .Q(g236), .D(g606), .test_si(n2162), 
        .test_so(n2161), .test_se(n2340) );
  dff_test_176 DFF_177 ( .CK(CK), .Q(g500), .D(g6292), .test_si(n2161), 
        .test_so(n2160), .test_se(n2341) );
  dff_test_177 DFF_178 ( .CK(CK), .Q(g205), .D(g5622), .test_si(n2160), 
        .test_so(n2159), .test_se(n2340) );
  dff_test_178 DFF_179 ( .CK(CK), .Q(g197), .D(g6287), .test_si(n2159), 
        .test_so(n2158), .test_se(n2341) );
  dff_test_179 DFF_180 ( .CK(CK), .Q(g666), .D(g4109), .test_si(n2158), 
        .test_so(n2157), .test_se(n2340) );
  dff_test_180 DFF_181 ( .CK(CK), .Q(g114), .D(g3727), .test_si(n2157), 
        .test_so(n2156), .test_se(n2341) );
  dff_test_181 DFF_182 ( .CK(CK), .Q(g524), .D(g6310), .test_si(n2156), 
        .test_so(n2155), .test_se(n2340) );
  dff_test_182 DFF_183 ( .CK(CK), .Q(g260), .D(g571), .test_si(n2155), 
        .test_so(n2154), .test_se(n2341) );
  dff_test_183 DFF_184 ( .CK(CK), .Q(g111), .D(g5701), .test_si(n2154), 
        .test_so(n2153), .test_se(n2340) );
  dff_test_184 DFF_185 ( .CK(CK), .Q(g131), .D(g4740), .test_si(n2153), 
        .test_so(n2152), .test_se(n2341) );
  dff_test_185 DFF_186 ( .CK(CK), .Q(g6688), .D(g6480), .test_si(n2152), 
        .test_so(n2151), .test_se(n2340) );
  dff_test_186 DFF_187 ( .CK(CK), .Q(g6691), .D(g6483), .test_si(n2151), 
        .test_so(n2150), .test_se(n2341) );
  dff_test_187 DFF_188 ( .CK(CK), .Q(g677), .D(g1), .test_si(n2150), .test_so(
        n2149), .test_se(n2340) );
  dff_test_188 DFF_189 ( .CK(CK), .Q(g582), .D(g6295), .test_si(n2149), 
        .test_so(n2148), .test_se(n2341) );
  dff_test_189 DFF_190 ( .CK(CK), .Q(g5468), .D(n656), .test_si(n2148), 
        .test_so(n2147), .test_se(n2340) );
  dff_test_190 DFF_191 ( .CK(CK), .Q(n2116), .D(n1247), .test_si(n2147), 
        .test_so(n2146), .test_se(n2341) );
  dff_test_191 DFF_192 ( .CK(CK), .Q(g193), .D(g5474), .test_si(n2146), 
        .test_so(n2145), .test_se(n2340) );
  dff_test_192 DFF_193 ( .CK(CK), .Q(g135), .D(g4752), .test_si(n2145), 
        .test_so(n2144), .test_se(n2341) );
  dff_test_193 DFF_194 ( .CK(CK), .Q(g382), .D(g5696), .test_si(n2144), 
        .test_so(n2143), .test_se(n2340) );
  dff_test_194 DFF_195 ( .CK(CK), .Q(g414), .D(g4447), .test_si(n2143), 
        .test_so(n2142), .test_se(n2341) );
  dff_test_195 DFF_196 ( .CK(CK), .Q(g434), .D(g4436), .test_si(n2142), 
        .test_so(n2141), .test_se(n2340) );
  dff_test_196 DFF_197 ( .CK(CK), .Q(g266), .D(g3910), .test_si(n2141), 
        .test_so(n2140), .test_se(n2341) );
  dff_test_197 DFF_198 ( .CK(CK), .Q(g49), .D(g6444), .test_si(n2140), 
        .test_so(n2139), .test_se(n2340) );
  dff_test_198 DFF_199 ( .CK(CK), .Q(g152), .D(g6109), .test_si(n2139), 
        .test_so(n2138), .test_se(n2341) );
  dff_test_199 DFF_200 ( .CK(CK), .Q(g692), .D(n1920), .test_si(n2138), 
        .test_so(n2137), .test_se(n2340) );
  dff_test_200 DFF_201 ( .CK(CK), .Q(g277), .D(g5625), .test_si(n2137), 
        .test_so(n2136), .test_se(n2341) );
  dff_test_201 DFF_202 ( .CK(CK), .Q(g127), .D(g6936), .test_si(n2136), 
        .test_so(n2135), .test_se(n2340) );
  dff_test_202 DFF_203 ( .CK(CK), .Q(g161), .D(g6113), .test_si(n2135), 
        .test_so(n2134), .test_se(n2341) );
  dff_test_203 DFF_204 ( .CK(CK), .Q(g512), .D(g6303), .test_si(n2134), 
        .test_so(n2133), .test_se(n2340) );
  dff_test_204 DFF_205 ( .CK(CK), .Q(g532), .D(g6301), .test_si(n2133), 
        .test_so(n2132), .test_se(n2341) );
  dff_test_205 DFF_206 ( .CK(CK), .Q(g64), .D(g6452), .test_si(n2132), 
        .test_so(n2131), .test_se(n2340) );
  dff_test_206 DFF_207 ( .CK(CK), .Q(g694), .D(g14), .test_si(n2131), 
        .test_so(n2130), .test_se(n2341) );
  dff_test_207 DFF_208 ( .CK(CK), .Q(g691), .D(n1915), .test_si(n2130), 
        .test_so(n2129), .test_se(n2340) );
  dff_test_208 DFF_209 ( .CK(CK), .Q(g1), .D(g6686), .test_si(n2129), 
        .test_so(n2128), .test_se(n2341) );
  dff_test_209 DFF_210 ( .CK(CK), .Q(g59), .D(g6450), .test_si(n2128), 
        .test_so(test_so), .test_se(n2340) );
  AO221X1 U1182 ( .IN1(n2022), .IN2(n1255), .IN3(g123), .IN4(n1256), .IN5(
        n1257), .Q(g6937) );
  OA22X1 U1186 ( .IN1(n1266), .IN2(n1155), .IN3(n1942), .IN4(n1910), .Q(n1263)
         );
  AO22X1 U1187 ( .IN1(n1269), .IN2(n2022), .IN3(n1270), .IN4(n1231), .Q(g6936)
         );
  AO22X1 U1188 ( .IN1(n1271), .IN2(n1209), .IN3(g127), .IN4(n1272), .Q(n1270)
         );
  NAND4X0 U1189 ( .IN1(g119), .IN2(n1273), .IN3(n1274), .IN4(n1233), .QN(n1272) );
  AO21X1 U1200 ( .IN1(n1966), .IN2(n1288), .IN3(n1290), .Q(n1280) );
  XNOR2X1 U1203 ( .IN1(n1051), .IN2(g284), .Q(n1297) );
  NAND3X0 U1204 ( .IN1(n1299), .IN2(n1300), .IN3(n1301), .QN(n1296) );
  XNOR2X1 U1205 ( .IN1(n1916), .IN2(g289), .Q(n1301) );
  NAND4X0 U1208 ( .IN1(n1302), .IN2(n1303), .IN3(n1304), .IN4(n1305), .QN(
        n1295) );
  XNOR2X1 U1209 ( .IN1(g680), .IN2(g286), .Q(n1305) );
  XNOR2X1 U1210 ( .IN1(g681), .IN2(g287), .Q(n1304) );
  XNOR2X1 U1211 ( .IN1(g684), .IN2(g290), .Q(n1303) );
  XNOR2X1 U1212 ( .IN1(g686), .IN2(g292), .Q(n1302) );
  AO222X1 U1217 ( .IN1(n1314), .IN2(g695), .IN3(n1315), .IN4(n1918), .IN5(
        n1909), .IN6(n1310), .Q(n1307) );
  OA22X1 U1218 ( .IN1(n1266), .IN2(n1168), .IN3(n2109), .IN4(n1962), .Q(n1279)
         );
  AO22X1 U1220 ( .IN1(n1319), .IN2(n2026), .IN3(n1320), .IN4(n1854), .Q(g6921)
         );
  AO21X1 U1221 ( .IN1(n1322), .IN2(g336), .IN3(n1240), .Q(n1320) );
  NAND4X0 U1223 ( .IN1(n1325), .IN2(n2053), .IN3(n1978), .IN4(n1242), .QN(
        n1324) );
  OR3X1 U1225 ( .IN1(n1753), .IN2(g332), .IN3(n1329), .Q(n1328) );
  AO221X1 U1227 ( .IN1(n1334), .IN2(n1335), .IN3(n1336), .IN4(n1337), .IN5(
        n2113), .Q(n1333) );
  AOI221X1 U1228 ( .IN1(n1336), .IN2(n1916), .IN3(n1334), .IN4(n1914), .IN5(
        n2089), .QN(n1339) );
  AO22X1 U1230 ( .IN1(n1950), .IN2(n2113), .IN3(n2090), .IN4(n1341), .Q(n1336)
         );
  OA22X1 U1231 ( .IN1(n1343), .IN2(n1342), .IN3(g337), .IN4(n1344), .Q(n1338)
         );
  OA221X1 U1232 ( .IN1(n1160), .IN2(n1960), .IN3(n1345), .IN4(n1346), .IN5(
        n2101), .Q(n1344) );
  OR2X1 U1233 ( .IN1(n1288), .IN2(n1171), .Q(n1346) );
  OA221X1 U1237 ( .IN1(n1192), .IN2(n1353), .IN3(n1108), .IN4(n1354), .IN5(
        n2087), .Q(n1352) );
  AOI221X1 U1238 ( .IN1(n1357), .IN2(n1916), .IN3(n1358), .IN4(n1914), .IN5(
        n2087), .QN(n1351) );
  OA221X1 U1239 ( .IN1(n1126), .IN2(n1353), .IN3(n1839), .IN4(n1354), .IN5(
        n2107), .Q(n1350) );
  AO22X1 U1240 ( .IN1(n2107), .IN2(n1051), .IN3(n2087), .IN4(n1359), .Q(n1354)
         );
  AO222X1 U1244 ( .IN1(n1798), .IN2(n1150), .IN3(n2087), .IN4(n1348), .IN5(
        g686), .IN6(n2106), .Q(n1362) );
  AO221X1 U1246 ( .IN1(n1358), .IN2(n1335), .IN3(n1337), .IN4(n1357), .IN5(
        n2106), .Q(n1361) );
  AO22X1 U1247 ( .IN1(n1950), .IN2(n2106), .IN3(n2088), .IN4(n1341), .Q(n1357)
         );
  AO22X1 U1250 ( .IN1(n2030), .IN2(n2108), .IN3(n1340), .IN4(n2088), .Q(n1358)
         );
  AO221X1 U1253 ( .IN1(n1363), .IN2(n1355), .IN3(n1364), .IN4(n1356), .IN5(
        n1960), .Q(n1331) );
  AO22X1 U1254 ( .IN1(g642), .IN2(n2085), .IN3(g230), .IN4(n2109), .Q(n1356)
         );
  AO22X1 U1255 ( .IN1(n1948), .IN2(n2043), .IN3(g218), .IN4(n2110), .Q(n1355)
         );
  AO221X1 U1256 ( .IN1(g679), .IN2(n1363), .IN3(g681), .IN4(n1364), .IN5(n2089), .Q(n1330) );
  AO22X1 U1257 ( .IN1(g680), .IN2(n2113), .IN3(n2091), .IN4(n1365), .Q(n1364)
         );
  AO22X1 U1259 ( .IN1(g678), .IN2(n2114), .IN3(n2090), .IN4(n1366), .Q(n1363)
         );
  NAND4X0 U1261 ( .IN1(n1971), .IN2(n1370), .IN3(n1369), .IN4(n1367), .QN(
        g6845) );
  OA221X1 U1262 ( .IN1(n1932), .IN2(n1899), .IN3(n1793), .IN4(n1837), .IN5(
        n1372), .Q(n1370) );
  AOI22X1 U1263 ( .IN1(n1788), .IN2(n1944), .IN3(g557), .IN4(n1972), .QN(n1372) );
  OA22X1 U1264 ( .IN1(n2103), .IN2(n1218), .IN3(n2104), .IN4(n1157), .Q(n1369)
         );
  NAND4X0 U1265 ( .IN1(n2073), .IN2(n1377), .IN3(n1376), .IN4(n1375), .QN(
        g6844) );
  OA221X1 U1266 ( .IN1(n1066), .IN2(n1835), .IN3(n1073), .IN4(n2101), .IN5(
        n1378), .Q(n1377) );
  AOI22X1 U1267 ( .IN1(n1788), .IN2(n1918), .IN3(g558), .IN4(n1972), .QN(n1378) );
  OA22X1 U1268 ( .IN1(n2102), .IN2(n1127), .IN3(n2105), .IN4(n1143), .Q(n1376)
         );
  AND2X1 U1278 ( .IN1(n1386), .IN2(n1146), .Q(n1385) );
  AOI21X1 U1286 ( .IN1(g211), .IN2(n1070), .IN3(n1399), .QN(n1392) );
  AO22X1 U1288 ( .IN1(n1386), .IN2(n1146), .IN3(n1401), .IN4(n1402), .Q(n1390)
         );
  XNOR2X1 U1289 ( .IN1(n1811), .IN2(n1099), .Q(n1401) );
  NAND4X0 U1291 ( .IN1(n1408), .IN2(n1407), .IN3(n1406), .IN4(n1409), .QN(
        n1405) );
  AOI22X1 U1295 ( .IN1(n1139), .IN2(n1410), .IN3(n1227), .IN4(n1414), .QN(
        n1413) );
  NAND3X0 U1298 ( .IN1(g211), .IN2(n1416), .IN3(g210), .QN(n1415) );
  NAND4X0 U1301 ( .IN1(n1424), .IN2(n1422), .IN3(n1423), .IN4(n1421), .QN(
        n1420) );
  AOI21X1 U1302 ( .IN1(n1169), .IN2(n1975), .IN3(n1140), .QN(n1424) );
  NAND4X0 U1305 ( .IN1(n1429), .IN2(n1140), .IN3(n1428), .IN4(n1427), .QN(
        n1419) );
  AOI22X1 U1306 ( .IN1(n1139), .IN2(n1426), .IN3(n1227), .IN4(n1975), .QN(
        n1429) );
  XOR2X1 U1309 ( .IN1(g471), .IN2(n1974), .Q(n1398) );
  NAND4X0 U1310 ( .IN1(n1971), .IN2(n1435), .IN3(n1434), .IN4(n1433), .QN(
        g6485) );
  OA221X1 U1311 ( .IN1(n1065), .IN2(n1932), .IN3(n1436), .IN4(n1793), .IN5(
        n1437), .Q(n1435) );
  OA22X1 U1313 ( .IN1(n2102), .IN2(n1163), .IN3(n2105), .IN4(n1197), .Q(n1434)
         );
  NAND4X0 U1314 ( .IN1(n2073), .IN2(n1440), .IN3(n1439), .IN4(n1438), .QN(
        g6483) );
  OA221X1 U1315 ( .IN1(n1063), .IN2(n1935), .IN3(n1096), .IN4(n2101), .IN5(
        n1441), .Q(n1440) );
  AOI22X1 U1316 ( .IN1(n1083), .IN2(n1909), .IN3(g560), .IN4(n1972), .QN(n1441) );
  OA22X1 U1317 ( .IN1(n2102), .IN2(n1170), .IN3(n2104), .IN4(n1153), .Q(n1439)
         );
  OA222X1 U1321 ( .IN1(n1895), .IN2(n1175), .IN3(n1149), .IN4(n1442), .IN5(
        n1155), .IN6(n1841), .Q(n1445) );
  AOI22X1 U1322 ( .IN1(n1084), .IN2(g554), .IN3(g561), .IN4(n1973), .QN(n1444)
         );
  AOI22X1 U1327 ( .IN1(n1084), .IN2(g551), .IN3(g562), .IN4(n1973), .QN(n1450)
         );
  NAND4X0 U1328 ( .IN1(n1457), .IN2(n1456), .IN3(n1455), .IN4(n1454), .QN(
        g6480) );
  OA222X1 U1330 ( .IN1(n1095), .IN2(n2100), .IN3(n2103), .IN4(n1151), .IN5(
        n2104), .IN6(n1203), .Q(n1456) );
  OA221X1 U1331 ( .IN1(n1987), .IN2(n1806), .IN3(n1797), .IN4(n1932), .IN5(
        n1461), .Q(n1455) );
  OA22X1 U1332 ( .IN1(n1961), .IN2(n1841), .IN3(n1895), .IN4(n1087), .Q(n1461)
         );
  AOI222X1 U1333 ( .IN1(g672), .IN2(n1050), .IN3(n1084), .IN4(g548), .IN5(g563), .IN6(n1973), .QN(n1454) );
  NAND4X0 U1334 ( .IN1(n1465), .IN2(n1464), .IN3(n1463), .IN4(n1462), .QN(
        g6479) );
  AND3X1 U1339 ( .IN1(n1473), .IN2(n1443), .IN3(n1448), .Q(n1472) );
  OA222X1 U1343 ( .IN1(n1094), .IN2(n2100), .IN3(n1869), .IN4(n1077), .IN5(
        n2105), .IN6(n1154), .Q(n1464) );
  NAND4X0 U1351 ( .IN1(n1481), .IN2(n1167), .IN3(n1993), .IN4(n1086), .QN(
        n1371) );
  AOI222X1 U1356 ( .IN1(n1050), .IN2(g669), .IN3(g545), .IN4(n1084), .IN5(
        n1973), .IN6(g564), .QN(n1462) );
  AND3X1 U1360 ( .IN1(n1479), .IN2(g683), .IN3(n1480), .Q(n1475) );
  NAND4X0 U1361 ( .IN1(n1868), .IN2(n1485), .IN3(g688), .IN4(n1486), .QN(n1471) );
  XNOR2X1 U1365 ( .IN1(n1088), .IN2(n1491), .Q(n1489) );
  AO21X1 U1367 ( .IN1(n2045), .IN2(n1497), .IN3(n2099), .Q(g6455) );
  AO21X1 U1374 ( .IN1(n1825), .IN2(n1508), .IN3(n1883), .Q(g6453) );
  AO221X1 U1376 ( .IN1(n1511), .IN2(n1120), .IN3(g386), .IN4(n1979), .IN5(
        n1507), .Q(n1510) );
  NOR3X0 U1377 ( .IN1(g59), .IN2(g64), .IN3(n1512), .QN(n1507) );
  AO21X1 U1378 ( .IN1(n1967), .IN2(n1514), .IN3(n2099), .Q(g6452) );
  OA222X1 U1380 ( .IN1(n2071), .IN2(n1216), .IN3(n1229), .IN4(n1861), .IN5(g59), .IN6(n1877), .Q(n1516) );
  AO21X1 U1381 ( .IN1(n1825), .IN2(n1517), .IN3(n2098), .Q(g6450) );
  AO21X1 U1391 ( .IN1(n2045), .IN2(n1529), .IN3(n2099), .Q(g6444) );
  XOR2X1 U1392 ( .IN1(g49), .IN2(n1530), .Q(n1529) );
  AO21X1 U1395 ( .IN1(n2045), .IN2(n1532), .IN3(n2098), .Q(g6440) );
  OA22X1 U1403 ( .IN1(n1844), .IN2(g84), .IN3(n1088), .IN4(n1496), .Q(n1540)
         );
  AND3X1 U1405 ( .IN1(n1521), .IN2(n1506), .IN3(g74), .Q(n1501) );
  AND3X1 U1406 ( .IN1(g49), .IN2(g361), .IN3(g54), .Q(n1521) );
  OA221X1 U1409 ( .IN1(n1326), .IN2(g314), .IN3(n1751), .IN4(n1857), .IN5(
        n1535), .Q(n1500) );
  AND4X1 U1410 ( .IN1(n1522), .IN2(n1229), .IN3(n1542), .IN4(n1226), .Q(n1502)
         );
  NOR3X0 U1411 ( .IN1(g49), .IN2(g54), .IN3(g361), .QN(n1522) );
  AO22X1 U1416 ( .IN1(n1792), .IN2(n1909), .IN3(n2095), .IN4(g516), .Q(g6307)
         );
  AO22X1 U1417 ( .IN1(n1792), .IN2(n1952), .IN3(g512), .IN4(n2097), .Q(g6303)
         );
  XNOR2X1 U1420 ( .IN1(g586), .IN2(n1549), .Q(n1552) );
  AO22X1 U1423 ( .IN1(n2016), .IN2(n1949), .IN3(g504), .IN4(n2095), .Q(g6296)
         );
  AO22X1 U1425 ( .IN1(g293), .IN2(n1856), .IN3(n1080), .IN4(n1951), .Q(g6294)
         );
  AND2X1 U1436 ( .IN1(g578), .IN2(n1562), .Q(n1555) );
  NAND4X0 U1441 ( .IN1(n1916), .IN2(n1212), .IN3(n1082), .IN4(n1566), .QN(
        n1551) );
  AND2X1 U1442 ( .IN1(n2025), .IN2(n1476), .Q(n1566) );
  NAND4X0 U1446 ( .IN1(n1476), .IN2(g677), .IN3(n1568), .IN4(n2025), .QN(n1550) );
  AND4X1 U1447 ( .IN1(n1485), .IN2(g684), .IN3(g685), .IN4(n1924), .Q(n1480)
         );
  OA221X1 U1450 ( .IN1(n1573), .IN2(n1165), .IN3(g586), .IN4(n1574), .IN5(
        n1575), .Q(n1572) );
  XNOR2X1 U1451 ( .IN1(g590), .IN2(g594), .Q(n1575) );
  OA22X1 U1452 ( .IN1(g582), .IN2(n1576), .IN3(n1577), .IN4(n1213), .Q(n1574)
         );
  OA22X1 U1453 ( .IN1(n1886), .IN2(n1903), .IN3(n1227), .IN4(n1196), .Q(n1577)
         );
  OA22X1 U1454 ( .IN1(n1886), .IN2(n1139), .IN3(n1177), .IN4(n1196), .Q(n1576)
         );
  OA22X1 U1455 ( .IN1(g582), .IN2(n1578), .IN3(n1579), .IN4(n1213), .Q(n1573)
         );
  OA22X1 U1456 ( .IN1(g578), .IN2(n1987), .IN3(n1169), .IN4(n1196), .Q(n1579)
         );
  NAND3X0 U1458 ( .IN1(g586), .IN2(g574), .IN3(g594), .QN(n1580) );
  OA22X1 U1461 ( .IN1(n1584), .IN2(n1057), .IN3(n2018), .IN4(n1214), .Q(n1583)
         );
  AO22X1 U1465 ( .IN1(g184), .IN2(n2017), .IN3(n1927), .IN4(n1591), .Q(n1589)
         );
  OA221X1 U1470 ( .IN1(g175), .IN2(n2018), .IN3(n2017), .IN4(n1598), .IN5(
        n1056), .Q(n1597) );
  XNOR3X1 U1475 ( .IN1(n1602), .IN2(n1603), .IN3(n1604), .Q(n1432) );
  XNOR3X1 U1476 ( .IN1(n1116), .IN2(g6688), .IN3(n1605), .Q(n1604) );
  XNOR2X1 U1477 ( .IN1(g6690), .IN2(g6691), .Q(n1605) );
  XNOR2X1 U1478 ( .IN1(n1166), .IN2(g6684), .Q(n1603) );
  XNOR2X1 U1479 ( .IN1(n1158), .IN2(g6686), .Q(n1602) );
  AND4X1 U1480 ( .IN1(g675), .IN2(n2082), .IN3(g676), .IN4(n1235), .Q(n1570)
         );
  AO22X1 U1482 ( .IN1(n1828), .IN2(g152), .IN3(n1608), .IN4(n1609), .Q(n1606)
         );
  OAI221X1 U1484 ( .IN1(n1138), .IN2(n2018), .IN3(n1610), .IN4(n1926), .IN5(
        n1220), .QN(n1608) );
  XNOR2X1 U1485 ( .IN1(g143), .IN2(n1954), .Q(n1610) );
  XNOR2X1 U1488 ( .IN1(n1185), .IN2(n1616), .Q(n1612) );
  AO21X1 U1489 ( .IN1(n1276), .IN2(n1234), .IN3(n2041), .Q(n1585) );
  AO221X1 U1490 ( .IN1(g398), .IN2(n1881), .IN3(g366), .IN4(n1988), .IN5(n2026), .Q(g5916) );
  OAI21X1 U1491 ( .IN1(n1619), .IN2(n1209), .IN3(n1620), .QN(g5701) );
  NAND4X0 U1492 ( .IN1(n1983), .IN2(n1230), .IN3(n1614), .IN4(n1209), .QN(
        n1620) );
  AO21X1 U1493 ( .IN1(n1983), .IN2(n1614), .IN3(n1820), .Q(n1617) );
  AOI21X1 U1494 ( .IN1(n1621), .IN2(n1615), .IN3(n1907), .QN(n1614) );
  AO21X1 U1495 ( .IN1(n1251), .IN2(n1867), .IN3(n1058), .Q(n1621) );
  AOI22X1 U1496 ( .IN1(n1919), .IN2(n1118), .IN3(g188), .IN4(n1874), .QN(n1613) );
  NAND4X0 U1497 ( .IN1(g179), .IN2(g170), .IN3(g161), .IN4(n1595), .QN(n1586)
         );
  AO22X1 U1505 ( .IN1(n1882), .IN2(g386), .IN3(n1807), .IN4(g390), .Q(g5698)
         );
  AO22X1 U1506 ( .IN1(n1882), .IN2(g382), .IN3(n1807), .IN4(g386), .Q(g5697)
         );
  AO22X1 U1507 ( .IN1(n1881), .IN2(g378), .IN3(n1807), .IN4(g382), .Q(g5696)
         );
  AO22X1 U1508 ( .IN1(n1882), .IN2(g374), .IN3(n1970), .IN4(g378), .Q(g5695)
         );
  AO22X1 U1509 ( .IN1(g370), .IN2(n1881), .IN3(n1970), .IN4(g374), .Q(g5694)
         );
  OA22X1 U1512 ( .IN1(n2091), .IN2(n1903), .IN3(n1623), .IN4(n1624), .Q(n1436)
         );
  AO22X1 U1514 ( .IN1(g695), .IN2(n2107), .IN3(n1628), .IN4(n1069), .Q(g5629)
         );
  NOR3X0 U1515 ( .IN1(n1630), .IN2(g209), .IN3(n1824), .QN(n1629) );
  AO22X1 U1516 ( .IN1(n1952), .IN2(n2114), .IN3(n1632), .IN4(n2090), .Q(g5628)
         );
  AO22X1 U1520 ( .IN1(n1952), .IN2(n2108), .IN3(n1637), .IN4(n2087), .Q(g5626)
         );
  AO22X1 U1522 ( .IN1(n1951), .IN2(n2107), .IN3(n1642), .IN4(n1641), .Q(g5624)
         );
  AO221X1 U1524 ( .IN1(n1105), .IN2(g193), .IN3(g148), .IN4(n1645), .IN5(n2022), .Q(g5583) );
  AO22X1 U1525 ( .IN1(n1909), .IN2(n1960), .IN3(n2091), .IN4(n1646), .Q(g5535)
         );
  AO22X1 U1528 ( .IN1(n1909), .IN2(n2107), .IN3(n2088), .IN4(n1648), .Q(g5533)
         );
  XNOR2X1 U1530 ( .IN1(n1631), .IN2(n1122), .Q(n1649) );
  AO22X1 U1531 ( .IN1(n2021), .IN2(n2114), .IN3(n1635), .IN4(n2028), .Q(g5532)
         );
  AND3X1 U1532 ( .IN1(n2090), .IN2(n1097), .IN3(n1801), .Q(n1635) );
  AND3X1 U1537 ( .IN1(n2088), .IN2(n1064), .IN3(n1069), .Q(n1642) );
  AO21X1 U1538 ( .IN1(n1974), .IN2(n1653), .IN3(n1070), .Q(n1639) );
  NOR3X0 U1540 ( .IN1(g211), .IN2(g471), .IN3(g210), .QN(n1653) );
  AO22X1 U1541 ( .IN1(n1105), .IN2(g184), .IN3(n1654), .IN4(g193), .Q(g5474)
         );
  AO22X1 U1542 ( .IN1(g175), .IN2(n1105), .IN3(n1654), .IN4(g184), .Q(g5473)
         );
  AO22X1 U1543 ( .IN1(n1105), .IN2(g166), .IN3(g175), .IN4(n1654), .Q(g5472)
         );
  AO22X1 U1544 ( .IN1(n1105), .IN2(g157), .IN3(n1654), .IN4(g166), .Q(g5471)
         );
  AO22X1 U1545 ( .IN1(g148), .IN2(n1105), .IN3(n1654), .IN4(g157), .Q(g5470)
         );
  AO21X1 U1547 ( .IN1(n1253), .IN2(n1235), .IN3(g669), .Q(g5386) );
  XNOR3X1 U1548 ( .IN1(n1655), .IN2(n1656), .IN3(n1930), .Q(n1253) );
  XOR2X1 U1549 ( .IN1(g4100), .IN2(g4099), .Q(n1656) );
  XOR3X1 U1550 ( .IN1(g4102), .IN2(g4101), .IN3(n1657), .Q(n1655) );
  XOR2X1 U1551 ( .IN1(g4105), .IN2(g4103), .Q(n1657) );
  AO21X1 U1553 ( .IN1(n1989), .IN2(n1180), .IN3(n1172), .Q(n1659) );
  AO221X1 U1554 ( .IN1(n1661), .IN2(n1135), .IN3(g349), .IN4(n1662), .IN5(
        n1131), .Q(g5295) );
  AO221X1 U1555 ( .IN1(n2077), .IN2(n1664), .IN3(n1135), .IN4(n1665), .IN5(
        n1131), .Q(g5291) );
  OR2X1 U1556 ( .IN1(n1665), .IN2(n1136), .Q(n1664) );
  NAND3X0 U1557 ( .IN1(n1945), .IN2(n1936), .IN3(n2077), .QN(n1665) );
  AO21X1 U1559 ( .IN1(n2078), .IN2(n1945), .IN3(n1936), .Q(n1667) );
  NAND3X0 U1569 ( .IN1(n1180), .IN2(n1172), .IN3(n1660), .QN(n1538) );
  NAND3X0 U1573 ( .IN1(n1176), .IN2(n1181), .IN3(g323), .QN(n1666) );
  AOI21X1 U1575 ( .IN1(n1800), .IN2(n1913), .IN3(g654), .QN(n1678) );
  AND3X1 U1579 ( .IN1(n1681), .IN2(g625), .IN3(g628), .Q(n1674) );
  AO21X1 U1582 ( .IN1(g139), .IN2(n1684), .IN3(n1104), .Q(g4757) );
  NAND3X0 U1585 ( .IN1(n1688), .IN2(n1103), .IN3(n1256), .QN(g4740) );
  XNOR2X1 U1588 ( .IN1(g625), .IN2(n1986), .Q(n1690) );
  AO22X1 U1593 ( .IN1(g426), .IN2(n2060), .IN3(n2064), .IN4(g422), .Q(g4458)
         );
  AO22X1 U1594 ( .IN1(g422), .IN2(n2057), .IN3(n1124), .IN4(g418), .Q(g4455)
         );
  AO22X1 U1595 ( .IN1(g445), .IN2(n2060), .IN3(n2064), .IN4(g449), .Q(g4454)
         );
  AO22X1 U1596 ( .IN1(g418), .IN2(n2058), .IN3(n2064), .IN4(g414), .Q(g4451)
         );
  AO22X1 U1597 ( .IN1(g449), .IN2(n2058), .IN3(n2062), .IN4(g453), .Q(g4450)
         );
  AO22X1 U1598 ( .IN1(g414), .IN2(n2058), .IN3(n2063), .IN4(g410), .Q(g4447)
         );
  AO22X1 U1599 ( .IN1(g453), .IN2(n2057), .IN3(n2061), .IN4(g457), .Q(g4446)
         );
  AO22X1 U1600 ( .IN1(g410), .IN2(n2059), .IN3(n2055), .IN4(g406), .Q(g4444)
         );
  AO22X1 U1601 ( .IN1(g457), .IN2(n2059), .IN3(n2063), .IN4(g461), .Q(g4443)
         );
  AO22X1 U1602 ( .IN1(g406), .IN2(n2115), .IN3(n2063), .IN4(g402), .Q(g4441)
         );
  AO22X1 U1603 ( .IN1(g461), .IN2(n2059), .IN3(n2063), .IN4(g430), .Q(g4440)
         );
  AO22X1 U1604 ( .IN1(g402), .IN2(n2059), .IN3(n1124), .IN4(n1698), .Q(g4438)
         );
  AO22X1 U1605 ( .IN1(g465), .IN2(n1811), .IN3(g471), .IN4(n1087), .Q(n1698)
         );
  AO22X1 U1606 ( .IN1(g434), .IN2(n2058), .IN3(n2062), .IN4(g437), .Q(g4436)
         );
  AO22X1 U1607 ( .IN1(g430), .IN2(n2060), .IN3(n2062), .IN4(g426), .Q(g4434)
         );
  AO22X1 U1608 ( .IN1(g437), .IN2(n2057), .IN3(n2061), .IN4(g441), .Q(g4433)
         );
  AO22X1 U1609 ( .IN1(g441), .IN2(n2060), .IN3(n2061), .IN4(g445), .Q(g4430)
         );
  NAND4X0 U1611 ( .IN1(n1700), .IN2(n1699), .IN3(n1701), .IN4(n1702), .QN(
        n1383) );
  XOR2X1 U1613 ( .IN1(g528), .IN2(g254), .Q(n1705) );
  XOR2X1 U1614 ( .IN1(g524), .IN2(g248), .Q(n1704) );
  XOR2X1 U1615 ( .IN1(g520), .IN2(g242), .Q(n1703) );
  NOR3X0 U1616 ( .IN1(n1708), .IN2(n1709), .IN3(n1707), .QN(n1701) );
  AND2X1 U1630 ( .IN1(g331), .IN2(n1691), .Q(g3731) );
  AND2X1 U1631 ( .IN1(n1691), .IN2(g328), .Q(g3730) );
  AND2X1 U1632 ( .IN1(g327), .IN2(n1691), .Q(g3729) );
  AND2X1 U1633 ( .IN1(g326), .IN2(n1691), .Q(g3728) );
  AND2X1 U1636 ( .IN1(g122), .IN2(n1694), .Q(g3727) );
  AND2X1 U1637 ( .IN1(n1694), .IN2(g119), .Q(g3726) );
  AND2X1 U1638 ( .IN1(g118), .IN2(n1694), .Q(g3725) );
  AND2X1 U1639 ( .IN1(g117), .IN2(n1694), .Q(g3724) );
  AOI21X1 U1641 ( .IN1(n1760), .IN2(n1252), .IN3(n1271), .QN(n1262) );
  OA22X1 U1643 ( .IN1(g3599), .IN2(n1110), .IN3(n1829), .IN4(n1190), .Q(n1718)
         );
  NOR3X0 U1645 ( .IN1(n1190), .IN2(n1310), .IN3(n1309), .QN(g2859) );
  AO22X1 U1646 ( .IN1(g2861), .IN2(n2039), .IN3(n1719), .IN4(g639), .Q(g2670)
         );
  OA22X1 U1647 ( .IN1(g489), .IN2(n1187), .IN3(g486), .IN4(n1111), .Q(g2433)
         );
  INVX0 U1650 ( .INP(1'b1), .ZN(g6728) );
  INVX0 U1652 ( .INP(1'b1), .ZN(g5692) );
  NAND3X2 U1654 ( .IN1(n1522), .IN2(n2071), .IN3(n2074), .QN(n1512) );
  DELLN1X2 U1655 ( .INP(n1535), .Z(n2075) );
  DELLN2X2 U1656 ( .INP(n1666), .Z(n2081) );
  DELLN1X2 U1657 ( .INP(n1550), .Z(n2096) );
  NOR2X1 U1658 ( .IN1(n1833), .IN2(n1516), .QN(n1515) );
  DELLN2X2 U1659 ( .INP(n1660), .Z(n1989) );
  INVX0 U1660 ( .INP(n2065), .ZN(n2067) );
  INVX0 U1661 ( .INP(n1643), .ZN(n1141) );
  DELLN1X2 U1662 ( .INP(n1176), .Z(n1945) );
  INVX0 U1663 ( .INP(n1813), .ZN(n1980) );
  NBUFFX2 U1664 ( .INP(n1550), .Z(n2097) );
  NBUFFX2 U1665 ( .INP(n1796), .Z(n2086) );
  XNOR2X2 U1666 ( .IN1(n1597), .IN2(n1188), .Q(n1596) );
  AO22X2 U1667 ( .IN1(g394), .IN2(n1882), .IN3(n1622), .IN4(g398), .Q(g5700)
         );
  DELLN2X2 U1668 ( .INP(n1410), .Z(n1816) );
  AO21X2 U1669 ( .IN1(n1541), .IN2(n1533), .IN3(n1538), .Q(n1537) );
  NAND3X4 U1670 ( .IN1(n1100), .IN2(n1890), .IN3(g465), .QN(n1559) );
  IBUFFX16 U1671 ( .INP(g276), .ZN(n2028) );
  AO22X2 U1672 ( .IN1(g551), .IN2(n1383), .IN3(n1851), .IN4(n1267), .Q(g6789)
         );
  AND2X1 U1673 ( .IN1(g279), .IN2(g278), .Q(n1878) );
  AND3X1 U1674 ( .IN1(n1938), .IN2(n1784), .IN3(n1487), .Q(n1925) );
  NBUFFX2 U1675 ( .INP(n1326), .Z(n2053) );
  AO22X1 U1676 ( .IN1(g606), .IN2(n2086), .IN3(g236), .IN4(n2111), .Q(n1341)
         );
  NAND3X0 U1677 ( .IN1(n1904), .IN2(n1243), .IN3(n1238), .QN(n1321) );
  INVX0 U1678 ( .INP(n2044), .ZN(n1894) );
  INVX0 U1679 ( .INP(n1762), .ZN(n1242) );
  NBUFFX2 U1680 ( .INP(g685), .Z(n1914) );
  NAND3X0 U1681 ( .IN1(n1086), .IN2(n1167), .IN3(n1993), .QN(n1345) );
  AO22X1 U1682 ( .IN1(n2030), .IN2(n1960), .IN3(n1340), .IN4(n2091), .Q(n1334)
         );
  XNOR2X1 U1683 ( .IN1(n1173), .IN2(g218), .Q(n1708) );
  XNOR2X1 U1684 ( .IN1(n1224), .IN2(g230), .Q(n1707) );
  XOR2X1 U1685 ( .IN1(g516), .IN2(g236), .Q(n1709) );
  NBUFFX2 U1686 ( .INP(n1374), .Z(n1840) );
  NAND3X1 U1687 ( .IN1(n1475), .IN2(g677), .IN3(n1476), .QN(n1443) );
  AO22X1 U1688 ( .IN1(n1760), .IN2(n2067), .IN3(n1262), .IN4(n1232), .Q(n1611)
         );
  OR2X1 U1689 ( .IN1(n1054), .IN2(n1904), .Q(n1541) );
  INVX0 U1690 ( .INP(n1801), .ZN(n1623) );
  DELLN1X2 U1691 ( .INP(g280), .Z(n1845) );
  AND3X1 U1692 ( .IN1(n1933), .IN2(n1997), .IN3(g279), .Q(n1957) );
  NBUFFX2 U1693 ( .INP(n1133), .Z(n1866) );
  INVX0 U1694 ( .INP(n1907), .ZN(n1259) );
  NBUFFX2 U1695 ( .INP(n1693), .Z(n2076) );
  AND2X1 U1696 ( .IN1(g582), .IN2(n1555), .Q(n1549) );
  AND3X1 U1697 ( .IN1(g654), .IN2(n1800), .IN3(n1679), .Q(n1676) );
  NBUFFX2 U1698 ( .INP(n1681), .Z(n1986) );
  OR2X1 U1699 ( .IN1(n2034), .IN2(n1992), .Q(n1631) );
  NBUFFX2 U1700 ( .INP(g128), .Z(n1870) );
  NBUFFX2 U1701 ( .INP(g114), .Z(n1871) );
  AO22X1 U1702 ( .IN1(n1951), .IN2(n2113), .IN3(n1635), .IN4(n1636), .Q(g5627)
         );
  AND2X1 U1703 ( .IN1(g702), .IN2(n2116), .Q(n1938) );
  NAND3X1 U1704 ( .IN1(n1205), .IN2(n1177), .IN3(n1940), .QN(n1428) );
  NAND3X0 U1705 ( .IN1(n1076), .IN2(n1199), .IN3(n1872), .QN(n1427) );
  NAND3X1 U1706 ( .IN1(n1205), .IN2(n1221), .IN3(n1940), .QN(n1421) );
  NAND3X0 U1707 ( .IN1(n1199), .IN2(n1228), .IN3(n1872), .QN(n1422) );
  NBUFFX2 U1708 ( .INP(n1796), .Z(n2085) );
  AO22X1 U1709 ( .IN1(n2108), .IN2(n1184), .IN3(n2088), .IN4(n1360), .Q(n1353)
         );
  OAI22X1 U1710 ( .IN1(n2109), .IN2(n1831), .IN3(g224), .IN4(n2044), .QN(n1360) );
  NAND3X0 U1711 ( .IN1(n1880), .IN2(n1177), .IN3(n1808), .QN(n1412) );
  NAND3X0 U1712 ( .IN1(n1880), .IN2(n1221), .IN3(n1808), .QN(n1406) );
  NAND3X0 U1713 ( .IN1(n2028), .IN2(n1228), .IN3(n1922), .QN(n1407) );
  AND2X1 U1714 ( .IN1(n1734), .IN2(n1430), .Q(n1838) );
  NAND3X1 U1715 ( .IN1(n1969), .IN2(n1212), .IN3(n1476), .QN(n1448) );
  NBUFFX2 U1716 ( .INP(g205), .Z(n1872) );
  AND3X1 U1717 ( .IN1(g691), .IN2(n1110), .IN3(g567), .Q(n2001) );
  XNOR2X1 U1718 ( .IN1(n1950), .IN2(g288), .Q(n1299) );
  XNOR2X1 U1719 ( .IN1(n1914), .IN2(g291), .Q(n1300) );
  XNOR2X1 U1720 ( .IN1(n1839), .IN2(g285), .Q(n1298) );
  NAND3X0 U1721 ( .IN1(n1798), .IN2(n1910), .IN3(n1082), .QN(n1288) );
  INVX0 U1722 ( .INP(g319), .ZN(n1244) );
  NBUFFX2 U1723 ( .INP(n1586), .Z(n1874) );
  NAND3X1 U1724 ( .IN1(n1868), .IN2(n1179), .IN3(n1480), .QN(n1449) );
  INVX0 U1725 ( .INP(g204), .ZN(n1199) );
  NBUFFX2 U1726 ( .INP(n1425), .Z(n1975) );
  NBUFFX2 U1727 ( .INP(n1480), .Z(n2025) );
  AO22X1 U1728 ( .IN1(g654), .IN2(n2085), .IN3(g254), .IN4(n2110), .Q(n1335)
         );
  AO22X1 U1729 ( .IN1(g646), .IN2(n2044), .IN3(g242), .IN4(n2110), .Q(n1337)
         );
  AO22X1 U1730 ( .IN1(n1948), .IN2(n2048), .IN3(g212), .IN4(n1894), .Q(n1366)
         );
  NOR2X0 U1731 ( .IN1(n1431), .IN2(n1152), .QN(n1399) );
  INVX0 U1732 ( .INP(g64), .ZN(n1226) );
  AND3X1 U1733 ( .IN1(g64), .IN2(g59), .IN3(g69), .Q(n1506) );
  AND3X1 U1734 ( .IN1(n2111), .IN2(n1787), .IN3(n1905), .Q(n1846) );
  AND3X1 U1735 ( .IN1(g680), .IN2(n1182), .IN3(n1051), .Q(n1486) );
  NAND3X0 U1736 ( .IN1(n1474), .IN2(n1182), .IN3(g678), .QN(n1458) );
  NAND3X0 U1737 ( .IN1(n1051), .IN2(n1182), .IN3(n1474), .QN(n1460) );
  INVX0 U1738 ( .INP(n1286), .ZN(n1048) );
  NAND3X0 U1739 ( .IN1(n1223), .IN2(n1188), .IN3(n1901), .QN(n1593) );
  NAND3X0 U1740 ( .IN1(g161), .IN2(n1855), .IN3(g170), .QN(n1592) );
  AND2X1 U1741 ( .IN1(g619), .IN2(n1712), .Q(n1696) );
  OA22X1 U1742 ( .IN1(n2106), .IN2(n1449), .IN3(n1225), .IN4(n1895), .Q(n1478)
         );
  INVX0 U1743 ( .INP(n1852), .ZN(n1869) );
  NBUFFX2 U1744 ( .INP(n1975), .Z(n1896) );
  INVX0 U1745 ( .INP(g69), .ZN(n1148) );
  NAND3X0 U1746 ( .IN1(n1082), .IN2(n1179), .IN3(n2025), .QN(n1553) );
  NAND3X0 U1747 ( .IN1(n1795), .IN2(n1243), .IN3(n2075), .QN(n1691) );
  INVX0 U1748 ( .INP(n1722), .ZN(n1237) );
  NOR2X0 U1749 ( .IN1(n1338), .IN2(n1339), .QN(n1332) );
  AOI22X1 U1750 ( .IN1(n1348), .IN2(n2091), .IN3(n1961), .IN4(g686), .QN(n1343) );
  NAND3X0 U1751 ( .IN1(n1259), .IN2(n1875), .IN3(g107), .QN(n1645) );
  NBUFFX2 U1752 ( .INP(n1545), .Z(n1985) );
  AND2X1 U1753 ( .IN1(n1717), .IN2(g616), .Q(n1712) );
  NBUFFX2 U1754 ( .INP(n1840), .Z(n2105) );
  NAND3X0 U1755 ( .IN1(n1889), .IN2(n1145), .IN3(n1626), .QN(n1625) );
  AND2X1 U1756 ( .IN1(n1618), .IN2(n1814), .Q(n1622) );
  INVX0 U1757 ( .INP(n2014), .ZN(n2016) );
  NBUFFX2 U1758 ( .INP(n1371), .Z(n1932) );
  AND2X1 U1759 ( .IN1(n1645), .IN2(n1231), .Q(n1654) );
  INVX0 U1760 ( .INP(n1611), .ZN(n1953) );
  NBUFFX2 U1761 ( .INP(n1512), .Z(n1877) );
  NBUFFX2 U1762 ( .INP(n1488), .Z(n1825) );
  NAND3X0 U1763 ( .IN1(n1791), .IN2(n1235), .IN3(g675), .QN(g6282) );
  NAND3X0 U1764 ( .IN1(n1801), .IN2(n1889), .IN3(n1647), .QN(n1646) );
  XNOR2X1 U1765 ( .IN1(n1845), .IN2(n1957), .Q(n1647) );
  INVX0 U1766 ( .INP(n1789), .ZN(g5531) );
  INVX0 U1767 ( .INP(n1797), .ZN(g5622) );
  DELLN1X2 U1768 ( .INP(g6), .Z(n1920) );
  NOR3X0 U1769 ( .IN1(n1751), .IN2(n1240), .IN3(n1329), .QN(n1382) );
  NAND3X0 U1770 ( .IN1(n1260), .IN2(n1261), .IN3(n1977), .QN(n1258) );
  XNOR2X1 U1771 ( .IN1(n1870), .IN2(n1871), .Q(n1682) );
  AO22X1 U1772 ( .IN1(g554), .IN2(n1383), .IN3(n1125), .IN4(n2023), .Q(g6790)
         );
  AO21X1 U1773 ( .IN1(n1398), .IN2(n1123), .IN3(n1394), .Q(n1416) );
  OA221X1 U1774 ( .IN1(n1373), .IN2(n1161), .IN3(n1897), .IN4(n1202), .IN5(
        n2072), .Q(n1453) );
  XNOR2X1 U1775 ( .IN1(n1109), .IN2(g606), .Q(n1710) );
  NOR3X0 U1776 ( .IN1(n1190), .IN2(n1913), .IN3(n1692), .QN(g4501) );
  XOR2X1 U1777 ( .IN1(n1892), .IN2(n1536), .Q(n1532) );
  NAND3X1 U1778 ( .IN1(n1069), .IN2(n1064), .IN3(n1649), .QN(n1648) );
  XOR2X1 U1779 ( .IN1(n1548), .IN2(g574), .Q(n1547) );
  INVX0 U1780 ( .INP(n1899), .ZN(g6792) );
  XNOR2X1 U1781 ( .IN1(n1676), .IN2(g571), .Q(n1675) );
  NAND3X0 U1782 ( .IN1(n1565), .IN2(n1178), .IN3(n1125), .QN(n1564) );
  OAI21X1 U1783 ( .IN1(n1809), .IN2(n1551), .IN3(n1556), .QN(g6293) );
  NAND3X0 U1784 ( .IN1(n1551), .IN2(n1557), .IN3(g536), .QN(n1556) );
  DELLN1X2 U1785 ( .INP(g24), .Z(n1912) );
  AO22X1 U1786 ( .IN1(g545), .IN2(n1383), .IN3(n1851), .IN4(n1941), .Q(g6787)
         );
  NAND3X0 U1787 ( .IN1(n1667), .IN2(n2081), .IN3(n1381), .QN(g5277) );
  NOR3X0 U1788 ( .IN1(n1249), .IN2(n1819), .IN3(n1680), .QN(g4872) );
  NAND3X0 U1789 ( .IN1(g283), .IN2(n1390), .IN3(g282), .QN(n1400) );
  NOR3X0 U1790 ( .IN1(n1902), .IN2(n1109), .IN3(n1713), .QN(g3844) );
  INVX0 U1791 ( .INP(n1962), .ZN(n655) );
  AO22X1 U1792 ( .IN1(n1882), .IN2(g390), .IN3(g394), .IN4(n1622), .Q(g5699)
         );
  AO22X1 U1793 ( .IN1(n1792), .IN2(n1951), .IN3(g508), .IN4(n2096), .Q(g6300)
         );
  AO22X1 U1794 ( .IN1(g548), .IN2(n1383), .IN3(n1851), .IN4(n1943), .Q(g6788)
         );
  AO22X1 U1795 ( .IN1(g366), .IN2(n1881), .IN3(g370), .IN4(n1622), .Q(g5693)
         );
  AO22X1 U1796 ( .IN1(n2015), .IN2(n2021), .IN3(g500), .IN4(n2097), .Q(g6292)
         );
  INVX0 U1797 ( .INP(n1942), .ZN(n656) );
  NOR3X0 U1798 ( .IN1(n1870), .IN2(g131), .IN3(n1215), .QN(n1687) );
  NBUFFX2 U1799 ( .INP(g2), .Z(n1915) );
  XNOR2X1 U1800 ( .IN1(n1800), .IN2(n1913), .Q(n1683) );
  NAND3X0 U1801 ( .IN1(n1178), .IN2(n1175), .IN3(n1125), .QN(n1697) );
  INVX0 U1802 ( .INP(n1947), .ZN(n1988) );
  INVX0 U1803 ( .INP(g688), .ZN(n1924) );
  NBUFFX2 U1804 ( .INP(n1924), .Z(n1993) );
  AND3X1 U1805 ( .IN1(n1891), .IN2(n2079), .IN3(n1534), .Q(n1883) );
  INVX0 U1806 ( .INP(n1697), .ZN(n2056) );
  AND2X1 U1807 ( .IN1(g586), .IN2(g574), .Q(n1727) );
  AND2X1 U1808 ( .IN1(n1239), .IN2(n1521), .Q(n1728) );
  AND2X1 U1809 ( .IN1(n1412), .IN2(n1091), .Q(n1729) );
  NAND3X0 U1810 ( .IN1(g679), .IN2(g678), .IN3(n1474), .QN(n1470) );
  AOI221X1 U1811 ( .IN1(n1280), .IN2(n1159), .IN3(n1281), .IN4(n1911), .IN5(
        n1803), .QN(n1730) );
  OR2X1 U1812 ( .IN1(g345), .IN2(g349), .Q(n1731) );
  OR2X1 U1813 ( .IN1(n1117), .IN2(n1119), .Q(n1732) );
  AND2X1 U1814 ( .IN1(n1445), .IN2(n1444), .Q(n1733) );
  AND2X1 U1815 ( .IN1(n1395), .IN2(g210), .Q(n1734) );
  AND2X1 U1816 ( .IN1(n1978), .IN2(g319), .Q(n1735) );
  AND3X1 U1817 ( .IN1(n1333), .IN2(n1331), .IN3(n1330), .Q(n1736) );
  AND2X1 U1818 ( .IN1(n1922), .IN2(n2028), .Q(n1737) );
  INVX0 U1819 ( .INP(n1997), .ZN(n1128) );
  INVX0 U1820 ( .INP(n1873), .ZN(n2064) );
  AND3X1 U1821 ( .IN1(n1086), .IN2(n1924), .IN3(n1167), .Q(n1738) );
  AND2X1 U1822 ( .IN1(n1501), .IN2(g79), .Q(n1739) );
  AND2X1 U1823 ( .IN1(n2069), .IN2(n1842), .Q(n1740) );
  AND3X1 U1824 ( .IN1(n1245), .IN2(n2116), .IN3(n1767), .Q(n1741) );
  AND2X1 U1825 ( .IN1(n2070), .IN2(n1537), .Q(n1833) );
  OR2X1 U1826 ( .IN1(n1555), .IN2(n1561), .Q(n1742) );
  NAND2X1 U1827 ( .IN1(n1815), .IN2(n1539), .QN(n1325) );
  OAI21X1 U1828 ( .IN1(n1243), .IN2(n1054), .IN3(n1328), .QN(n1743) );
  AND3X1 U1829 ( .IN1(n1237), .IN2(g328), .IN3(n1324), .Q(n1744) );
  OR2X1 U1830 ( .IN1(n1220), .IN2(n1185), .Q(n1745) );
  AND2X1 U1831 ( .IN1(g682), .IN2(g677), .Q(n1746) );
  OAI21X1 U1832 ( .IN1(n1537), .IN2(n1540), .IN3(n1854), .QN(n1747) );
  NAND2X0 U1833 ( .IN1(n1795), .IN2(n1740), .QN(n1535) );
  NBUFFX2 U1834 ( .INP(n1752), .Z(n2052) );
  INVX0 U1835 ( .INP(n1747), .ZN(n1488) );
  INVX0 U1836 ( .INP(n1747), .ZN(n2045) );
  NAND2X0 U1837 ( .IN1(n1523), .IN2(n1967), .QN(n1748) );
  INVX0 U1838 ( .INP(n1883), .ZN(n1749) );
  NAND2X0 U1839 ( .IN1(n1748), .IN2(n1749), .QN(g6447) );
  XNOR2X1 U1840 ( .IN1(n1524), .IN2(g54), .Q(n1523) );
  INVX0 U1841 ( .INP(n1843), .ZN(n1968) );
  NAND2X0 U1842 ( .IN1(n2045), .IN2(n1489), .QN(n1750) );
  NAND2X0 U1843 ( .IN1(n1750), .IN2(n1749), .QN(g6456) );
  NBUFFX2 U1844 ( .INP(n2052), .Z(n1751) );
  NBUFFX2 U1845 ( .INP(g306), .Z(n1752) );
  INVX0 U1846 ( .INP(n1978), .ZN(n1753) );
  NBUFFX2 U1847 ( .INP(n2070), .Z(n1754) );
  NBUFFX2 U1848 ( .INP(n1238), .Z(n1978) );
  NAND2X0 U1849 ( .IN1(n1503), .IN2(n1967), .QN(n1755) );
  INVX0 U1850 ( .INP(n2098), .ZN(n1756) );
  NAND2X0 U1851 ( .IN1(n1755), .IN2(n1756), .QN(g6454) );
  INVX0 U1852 ( .INP(g314), .ZN(n1243) );
  AND3X1 U1853 ( .IN1(n1892), .IN2(n1968), .IN3(g49), .Q(n1999) );
  NAND3X0 U1854 ( .IN1(n2050), .IN2(n1244), .IN3(g301), .QN(n1533) );
  INVX0 U1855 ( .INP(g46), .ZN(n1757) );
  INVX0 U1856 ( .INP(n1757), .ZN(g4109) );
  INVX0 U1857 ( .INP(g94), .ZN(n1759) );
  INVX0 U1858 ( .INP(n1759), .ZN(n1760) );
  INVX0 U1859 ( .INP(g310), .ZN(n1761) );
  INVX0 U1860 ( .INP(n1761), .ZN(n1762) );
  INVX0 U1861 ( .INP(g102), .ZN(n1232) );
  INVX0 U1862 ( .INP(g45), .ZN(n1763) );
  INVX0 U1863 ( .INP(n1763), .ZN(g4108) );
  INVX0 U1864 ( .INP(n1252), .ZN(n1765) );
  INVX0 U1865 ( .INP(g702), .ZN(n1766) );
  INVX0 U1866 ( .INP(n1766), .ZN(n1767) );
  INVX0 U1867 ( .INP(g42), .ZN(n1768) );
  INVX0 U1868 ( .INP(n1768), .ZN(g4106) );
  INVX0 U1869 ( .INP(g40), .ZN(n1770) );
  INVX0 U1870 ( .INP(n1770), .ZN(g4105) );
  INVX0 U1871 ( .INP(g39), .ZN(n1772) );
  INVX0 U1872 ( .INP(n1772), .ZN(g4103) );
  INVX0 U1873 ( .INP(g38), .ZN(n1774) );
  INVX0 U1874 ( .INP(n1774), .ZN(g4102) );
  INVX0 U1875 ( .INP(g37), .ZN(n1776) );
  INVX0 U1876 ( .INP(n1776), .ZN(g4101) );
  INVX0 U1877 ( .INP(g36), .ZN(n1778) );
  INVX0 U1878 ( .INP(n1778), .ZN(g4100) );
  INVX0 U1879 ( .INP(g32), .ZN(n1780) );
  INVX0 U1880 ( .INP(n1780), .ZN(g4099) );
  INVX0 U1881 ( .INP(g41), .ZN(n1782) );
  INVX0 U1882 ( .INP(n1782), .ZN(n1783) );
  INVX0 U1883 ( .INP(n1782), .ZN(n1784) );
  AND3X1 U1884 ( .IN1(n1185), .IN2(n1220), .IN3(n1611), .Q(n1594) );
  XNOR2X2 U1885 ( .IN1(g18), .IN2(g14), .Q(n1671) );
  AO21X1 U1886 ( .IN1(n1290), .IN2(n1482), .IN3(n1931), .Q(n1442) );
  AO21X1 U1887 ( .IN1(n1290), .IN2(n1482), .IN3(n1931), .Q(n1806) );
  OA221X1 U1888 ( .IN1(n2103), .IN2(n1142), .IN3(n1897), .IN4(n1224), .IN5(
        n2072), .Q(n1447) );
  OA222X1 U1889 ( .IN1(n1059), .IN2(n1835), .IN3(n2105), .IN4(n1217), .IN5(
        n1092), .IN6(n2100), .Q(n1446) );
  INVX0 U1890 ( .INP(n1939), .ZN(n1940) );
  NAND2X1 U1891 ( .IN1(n1391), .IN2(g210), .QN(n1785) );
  NAND2X0 U1892 ( .IN1(n1392), .IN2(g211), .QN(n1786) );
  NAND3X0 U1893 ( .IN1(n1785), .IN2(n1786), .IN3(n1393), .QN(n1316) );
  AND2X1 U1894 ( .IN1(n1484), .IN2(g662), .Q(n1787) );
  INVX0 U1895 ( .INP(n1806), .ZN(n1788) );
  INVX0 U1896 ( .INP(n1651), .ZN(n1099) );
  AOI22X2 U1897 ( .IN1(n2021), .IN2(n2108), .IN3(n1642), .IN4(n1199), .QN(
        n1789) );
  XNOR3X1 U1898 ( .IN1(n1826), .IN2(g48), .IN3(n1790), .Q(n1569) );
  XOR3X1 U1899 ( .IN1(g10), .IN2(g1), .IN3(n1671), .Q(n1790) );
  NAND2X0 U1900 ( .IN1(n1846), .IN2(n1847), .QN(n1347) );
  DELLN1X2 U1901 ( .INP(n1905), .Z(n1791) );
  INVX0 U1902 ( .INP(n1935), .ZN(n1834) );
  NBUFFX2 U1903 ( .INP(n1079), .Z(n1792) );
  NAND2X0 U1904 ( .IN1(n1846), .IN2(n1847), .QN(n1793) );
  AO221X1 U1905 ( .IN1(n1610), .IN2(n2018), .IN3(n1106), .IN4(n1138), .IN5(
        n1220), .Q(n1609) );
  NBUFFX2 U1906 ( .INP(g197), .Z(n1794) );
  NAND3X0 U1907 ( .IN1(n2067), .IN2(n1234), .IN3(n1876), .QN(n1615) );
  NAND2X0 U1908 ( .IN1(n1813), .IN2(n1728), .QN(n1513) );
  NBUFFX2 U1909 ( .INP(n1241), .Z(n1795) );
  NBUFFX2 U1910 ( .INP(g658), .Z(n1796) );
  AOI22X1 U1911 ( .IN1(n1949), .IN2(n2108), .IN3(n1644), .IN4(n1642), .QN(
        n1797) );
  XNOR2X1 U1912 ( .IN1(n1504), .IN2(g74), .Q(n1503) );
  NBUFFX2 U1913 ( .INP(n1814), .Z(n1854) );
  INVX0 U1914 ( .INP(n1160), .ZN(n1798) );
  INVX0 U1915 ( .INP(g662), .ZN(n1160) );
  NAND2X0 U1916 ( .IN1(n2030), .IN2(n1159), .QN(n1823) );
  AOI22X1 U1917 ( .IN1(n1083), .IN2(n1810), .IN3(g559), .IN4(n1972), .QN(n1437) );
  INVX0 U1918 ( .INP(g650), .ZN(n1799) );
  INVX0 U1919 ( .INP(n1799), .ZN(n1800) );
  AND2X1 U1920 ( .IN1(n2048), .IN2(g598), .Q(n1309) );
  NBUFFX2 U1921 ( .INP(g697), .Z(n1944) );
  NOR2X0 U1922 ( .IN1(n1388), .IN2(n1802), .QN(n1801) );
  NOR4X0 U1923 ( .IN1(n1994), .IN2(g282), .IN3(g283), .IN4(g478), .QN(n1802)
         );
  AO22X1 U1924 ( .IN1(n1048), .IN2(n1283), .IN3(n1284), .IN4(n2086), .Q(n1803)
         );
  AND2X1 U1925 ( .IN1(n1787), .IN2(n2111), .Q(n1804) );
  NBUFFX2 U1926 ( .INP(n1500), .Z(n1843) );
  INVX0 U1927 ( .INP(n1651), .ZN(n1994) );
  AND2X1 U1928 ( .IN1(n1471), .IN2(n1470), .Q(n1805) );
  AND3X1 U1929 ( .IN1(n1934), .IN2(n1347), .IN3(n1805), .Q(n1469) );
  INVX0 U1930 ( .INP(n1998), .ZN(n2071) );
  NOR3X0 U1931 ( .IN1(g361), .IN2(g49), .IN3(n1968), .QN(n2000) );
  NAND2X1 U1932 ( .IN1(n1510), .IN2(n2080), .QN(n1509) );
  AND3X1 U1933 ( .IN1(g682), .IN2(n1212), .IN3(n1969), .Q(n1852) );
  AO22X1 U1934 ( .IN1(n1918), .IN2(n2108), .IN3(n1941), .IN4(n2088), .Q(g6791)
         );
  NBUFFX2 U1935 ( .INP(n1622), .Z(n1807) );
  INVX0 U1936 ( .INP(n1754), .ZN(n1981) );
  NBUFFX2 U1937 ( .INP(n1929), .Z(n1808) );
  NBUFFX2 U1938 ( .INP(n1200), .Z(n2111) );
  NBUFFX2 U1939 ( .INP(n1200), .Z(n2109) );
  AND2X1 U1940 ( .IN1(g687), .IN2(n1738), .Q(n1847) );
  INVX0 U1941 ( .INP(n1951), .ZN(n1809) );
  NBUFFX2 U1942 ( .INP(g692), .Z(n1951) );
  INVX0 U1943 ( .INP(n1903), .ZN(n1810) );
  NBUFFX2 U1944 ( .INP(n1076), .Z(n1903) );
  XNOR2X2 U1945 ( .IN1(g281), .IN2(n1193), .Q(n1402) );
  NBUFFX2 U1946 ( .INP(g478), .Z(n1811) );
  AND2X1 U1947 ( .IN1(n1309), .IN2(g634), .Q(n1306) );
  AND3X1 U1948 ( .IN1(n1374), .IN2(n1373), .IN3(n1371), .Q(n1812) );
  AND2X1 U1949 ( .IN1(n1469), .IN2(n1812), .Q(n1468) );
  INVX0 U1950 ( .INP(n1858), .ZN(n1813) );
  INVX0 U1951 ( .INP(n2071), .ZN(n1858) );
  AND3X1 U1952 ( .IN1(g1293), .IN2(n2082), .IN3(n1767), .Q(n1484) );
  NBUFFX2 U1953 ( .INP(n1500), .Z(n2074) );
  NAND2X1 U1954 ( .IN1(n1505), .IN2(n2080), .QN(n1504) );
  NAND2X1 U1955 ( .IN1(n1884), .IN2(n1525), .QN(n1524) );
  NBUFFX2 U1956 ( .INP(n1321), .Z(n1814) );
  NBUFFX2 U1957 ( .INP(n1840), .Z(n2104) );
  AND2X1 U1958 ( .IN1(n1238), .IN2(n1244), .Q(n1815) );
  NAND3X1 U1959 ( .IN1(n1520), .IN2(n1877), .IN3(n1861), .QN(n1519) );
  AO222X1 U1960 ( .IN1(n2026), .IN2(n1379), .IN3(n1380), .IN4(n1866), .IN5(
        n1381), .IN6(g332), .Q(g6795) );
  OA221X1 U1961 ( .IN1(g370), .IN2(n1754), .IN3(n1980), .IN4(n1531), .IN5(
        n1494), .Q(n1530) );
  OA221X1 U1962 ( .IN1(g398), .IN2(n1859), .IN3(n1980), .IN4(n1493), .IN5(
        n1494), .Q(n1491) );
  NBUFFX2 U1963 ( .INP(n1070), .Z(n1817) );
  INVX0 U1964 ( .INP(n1817), .ZN(n1818) );
  AO22X1 U1965 ( .IN1(g650), .IN2(n2085), .IN3(g248), .IN4(n2109), .Q(n1340)
         );
  NAND2X0 U1966 ( .IN1(n1076), .IN2(n1737), .QN(n1411) );
  NBUFFX2 U1967 ( .INP(g277), .Z(n1922) );
  NBUFFX2 U1968 ( .INP(n1674), .Z(n1819) );
  NBUFFX2 U1969 ( .INP(n1254), .Z(n1820) );
  INVX0 U1970 ( .INP(n1852), .ZN(n1373) );
  AOI22X1 U1971 ( .IN1(n1944), .IN2(n2114), .IN3(n1268), .IN4(n2091), .QN(
        n1821) );
  IBUFFX16 U1972 ( .INP(n1821), .ZN(g6794) );
  NAND2X0 U1973 ( .IN1(n1279), .IN2(n1264), .QN(n1822) );
  NAND3X0 U1974 ( .IN1(n1822), .IN2(n1823), .IN3(n1730), .QN(n1269) );
  NBUFFX2 U1975 ( .INP(n1399), .Z(n1824) );
  AO22X1 U1976 ( .IN1(n1817), .IN2(n1087), .IN3(g465), .IN4(n1850), .Q(n1565)
         );
  NAND2X0 U1977 ( .IN1(n1239), .IN2(n1739), .QN(n1496) );
  XOR3X1 U1978 ( .IN1(g24), .IN2(g2), .IN3(n1672), .Q(n1826) );
  NAND2X0 U1979 ( .IN1(n1905), .IN2(n1804), .QN(n1865) );
  XOR2X1 U1980 ( .IN1(n1515), .IN2(g64), .Q(n1514) );
  AND2X1 U1981 ( .IN1(g622), .IN2(g619), .Q(n1827) );
  NAND2X1 U1982 ( .IN1(n1519), .IN2(n1884), .QN(n1518) );
  INVX0 U1983 ( .INP(n2084), .ZN(n1200) );
  INVX0 U1984 ( .INP(n1056), .ZN(n1828) );
  INVX0 U1985 ( .INP(n1607), .ZN(n1056) );
  INVX0 U1986 ( .INP(g634), .ZN(n1829) );
  INVX0 U1987 ( .INP(n1829), .ZN(n1830) );
  INVX0 U1988 ( .INP(n1829), .ZN(n1831) );
  NBUFFX2 U1989 ( .INP(n1316), .Z(n1943) );
  INVX0 U1990 ( .INP(n1824), .ZN(n1064) );
  AND2X1 U1991 ( .IN1(n1397), .IN2(g210), .Q(n1832) );
  IBUFFX16 U1992 ( .INP(n1998), .ZN(n2070) );
  NAND2X1 U1993 ( .IN1(n1832), .IN2(n1393), .QN(n1396) );
  NAND2X0 U1994 ( .IN1(n1332), .IN2(n1736), .QN(n1319) );
  NAND3X0 U1995 ( .IN1(n1261), .IN2(n1232), .IN3(n1977), .QN(n1694) );
  NBUFFX2 U1996 ( .INP(n1262), .Z(n1977) );
  NAND3X0 U1997 ( .IN1(n1447), .IN2(n1733), .IN3(n1446), .QN(g6482) );
  NOR2X0 U1998 ( .IN1(n1693), .IN2(n1732), .QN(n1679) );
  INVX0 U1999 ( .INP(n1834), .ZN(n1835) );
  AND2X1 U2000 ( .IN1(n1874), .IN2(n1919), .Q(n1584) );
  AND2X1 U2001 ( .IN1(n1502), .IN2(n1195), .Q(n1836) );
  INVX0 U2002 ( .INP(g6794), .ZN(n1837) );
  NBUFFX2 U2003 ( .INP(n1268), .Z(n2023) );
  XNOR2X2 U2004 ( .IN1(g209), .IN2(g208), .Q(n1430) );
  NBUFFX2 U2005 ( .INP(n1182), .Z(n1839) );
  INVX0 U2006 ( .INP(n1652), .ZN(n1100) );
  NBUFFX2 U2007 ( .INP(n1449), .Z(n1841) );
  INVX0 U2008 ( .INP(n1761), .ZN(n1842) );
  NAND2X0 U2009 ( .IN1(n2074), .IN2(n1836), .QN(n1844) );
  OAI21X1 U2010 ( .IN1(n1537), .IN2(n1540), .IN3(n1854), .QN(n2079) );
  INVX0 U2011 ( .INP(n1843), .ZN(n1239) );
  NAND2X0 U2012 ( .IN1(n1969), .IN2(n1746), .QN(n1374) );
  NAND2X1 U2013 ( .IN1(n1263), .IN2(n1264), .QN(n1955) );
  NAND2X1 U2014 ( .IN1(g282), .IN2(n1384), .QN(n1848) );
  NAND2X0 U2015 ( .IN1(g283), .IN2(n1101), .QN(n1849) );
  NAND2X1 U2016 ( .IN1(n1848), .IN2(n1849), .QN(n1268) );
  DELLN1X2 U2017 ( .INP(n1388), .Z(n1850) );
  NOR2X0 U2018 ( .IN1(n1652), .IN2(n1890), .QN(n1388) );
  AO22X2 U2019 ( .IN1(n1918), .IN2(n1961), .IN3(n2090), .IN4(n1267), .Q(g6793)
         );
  NAND2X1 U2020 ( .IN1(n1405), .IN2(n1404), .QN(n1403) );
  NBUFFX2 U2021 ( .INP(n1125), .Z(n1851) );
  XNOR2X1 U2022 ( .IN1(n1225), .IN2(g260), .Q(n1706) );
  INVX0 U2023 ( .INP(n1389), .ZN(n1889) );
  INVX0 U2024 ( .INP(g89), .ZN(n1875) );
  NAND3X0 U2025 ( .IN1(n1413), .IN2(n1729), .IN3(n1411), .QN(n1404) );
  AND2X1 U2026 ( .IN1(n1853), .IN2(n1430), .Q(n1394) );
  XOR2X1 U2027 ( .IN1(n1418), .IN2(g471), .Q(n1853) );
  NAND2X0 U2028 ( .IN1(n1159), .IN2(n1121), .QN(n1956) );
  AOI21X1 U2029 ( .IN1(n1997), .IN2(n1933), .IN3(g279), .QN(n1634) );
  NAND2X1 U2030 ( .IN1(n1387), .IN2(g282), .QN(n1887) );
  NBUFFX2 U2031 ( .INP(n1595), .Z(n1855) );
  NAND2X0 U2032 ( .IN1(n1741), .IN2(n1483), .QN(n1567) );
  NBUFFX2 U2033 ( .INP(n1553), .Z(n1856) );
  AO221X1 U2034 ( .IN1(n1287), .IN2(n1126), .IN3(n1283), .IN4(n1839), .IN5(
        n1189), .Q(n1281) );
  AO22X1 U2035 ( .IN1(g571), .IN2(n1796), .IN3(g260), .IN4(n1911), .Q(n1348)
         );
  AO22X1 U2036 ( .IN1(n2085), .IN2(n1830), .IN3(g224), .IN4(n1910), .Q(n1365)
         );
  NAND2X1 U2037 ( .IN1(g281), .IN2(n1627), .QN(n1652) );
  NBUFFX2 U2038 ( .INP(n2069), .Z(n1857) );
  OA221X1 U2039 ( .IN1(g394), .IN2(n1859), .IN3(n1981), .IN4(n1499), .IN5(
        n1494), .Q(n1991) );
  OA22X1 U2040 ( .IN1(n2074), .IN2(n1501), .IN3(n1968), .IN4(n1502), .Q(n1499)
         );
  XNOR2X1 U2041 ( .IN1(n1892), .IN2(n1968), .Q(n1531) );
  XOR2X1 U2042 ( .IN1(n1518), .IN2(n1229), .Q(n1517) );
  INVX0 U2043 ( .INP(n1858), .ZN(n1859) );
  INVX0 U2044 ( .INP(n1513), .ZN(n1860) );
  INVX0 U2045 ( .INP(n1860), .ZN(n1861) );
  AND2X1 U2046 ( .IN1(n2038), .IN2(g610), .Q(n1862) );
  AND2X1 U2047 ( .IN1(n1862), .IN2(n1863), .Q(n1681) );
  AND2X1 U2048 ( .IN1(n1827), .IN2(g616), .Q(n1863) );
  XOR2X1 U2049 ( .IN1(n1509), .IN2(n1148), .Q(n1508) );
  XOR2X1 U2050 ( .IN1(g224), .IN2(n1202), .Q(n1700) );
  DELLN1X2 U2051 ( .INP(g689), .Z(n1928) );
  XOR2X1 U2052 ( .IN1(g212), .IN2(n1204), .Q(n1699) );
  AO22X1 U2053 ( .IN1(g254), .IN2(g248), .IN3(g242), .IN4(g236), .Q(n1318) );
  AOI222X1 U2054 ( .IN1(n1944), .IN2(n1306), .IN3(n1831), .IN4(n1307), .IN5(
        n1308), .IN6(n1829), .QN(n1293) );
  AO22X1 U2055 ( .IN1(g297), .IN2(n1553), .IN3(n1080), .IN4(n1952), .Q(g6298)
         );
  AO22X1 U2056 ( .IN1(n2090), .IN2(n1856), .IN3(n1080), .IN4(n1949), .Q(g6290)
         );
  AND2X1 U2057 ( .IN1(n1700), .IN2(n1699), .Q(n1864) );
  OA222X1 U2058 ( .IN1(n1062), .IN2(n1835), .IN3(n2104), .IN4(n1156), .IN5(
        n1093), .IN6(n2100), .Q(n1452) );
  INVX0 U2059 ( .INP(n1765), .ZN(n1867) );
  NBUFFX2 U2060 ( .INP(n1925), .Z(n1868) );
  NBUFFX2 U2061 ( .INP(n1483), .Z(n1905) );
  XNOR2X1 U2062 ( .IN1(n1101), .IN2(n1385), .Q(n1384) );
  OAI22X1 U2063 ( .IN1(n2110), .IN2(g567), .IN3(g212), .IN4(n2085), .QN(n1359)
         );
  INVX0 U2064 ( .INP(n2056), .ZN(n1873) );
  NOR2X0 U2065 ( .IN1(n1611), .IN2(n1745), .QN(n1595) );
  INVX0 U2066 ( .INP(n1250), .ZN(n1876) );
  OAI21X1 U2067 ( .IN1(n1234), .IN2(n2024), .IN3(n2066), .QN(n1275) );
  AND2X1 U2068 ( .IN1(n1414), .IN2(n1878), .Q(n1627) );
  IBUFFX16 U2069 ( .INP(n1222), .ZN(n1879) );
  INVX0 U2070 ( .INP(n1879), .ZN(n1880) );
  DELLN1X2 U2071 ( .INP(n1276), .Z(n2024) );
  INVX0 U2072 ( .INP(n1988), .ZN(n1881) );
  INVX0 U2073 ( .INP(n1988), .ZN(n1882) );
  XOR2X1 U2074 ( .IN1(n1223), .IN2(n1600), .Q(n1599) );
  XOR2X1 U2075 ( .IN1(n1118), .IN2(n1583), .Q(n1581) );
  XOR2X1 U2076 ( .IN1(n1589), .IN2(g179), .Q(n1588) );
  AND4X1 U2077 ( .IN1(g688), .IN2(n1925), .IN3(n1485), .IN4(n1184), .Q(n1474)
         );
  INVX0 U2078 ( .INP(n1833), .ZN(n1884) );
  NBUFFX2 U2079 ( .INP(n1551), .Z(n1885) );
  XOR2X1 U2080 ( .IN1(g6), .IN2(g28), .Q(n1672) );
  INVX0 U2081 ( .INP(n1585), .ZN(n1106) );
  NAND2X1 U2082 ( .IN1(n2070), .IN2(n1537), .QN(n1494) );
  INVX0 U2083 ( .INP(n1196), .ZN(n1886) );
  INVX0 U2084 ( .INP(g578), .ZN(n1196) );
  NAND2X0 U2085 ( .IN1(n1850), .IN2(g283), .QN(n1888) );
  NAND3X0 U2086 ( .IN1(n1887), .IN2(n1888), .IN3(n1097), .QN(n1267) );
  INVX0 U2087 ( .INP(g280), .ZN(n1890) );
  NOR4X0 U2088 ( .IN1(n1995), .IN2(g282), .IN3(g283), .IN4(n1811), .QN(n1389)
         );
  AND2X1 U2089 ( .IN1(n2053), .IN2(n1533), .Q(n1891) );
  AND3X1 U2090 ( .IN1(n1534), .IN2(n1891), .IN3(n2079), .Q(n1490) );
  NBUFFX2 U2091 ( .INP(g361), .Z(n1892) );
  AND2X1 U2092 ( .IN1(n1613), .IN2(n2068), .Q(n1893) );
  INVX0 U2093 ( .INP(n1906), .ZN(n2054) );
  NBUFFX2 U2094 ( .INP(n1448), .Z(n1895) );
  NOR2X0 U2095 ( .IN1(n1643), .IN2(n2035), .QN(n1560) );
  NBUFFX2 U2096 ( .INP(n1443), .Z(n1897) );
  AOI221X1 U2097 ( .IN1(n1280), .IN2(n1159), .IN3(n1281), .IN4(n1911), .IN5(
        n1282), .QN(n1898) );
  NAND2X1 U2098 ( .IN1(n1420), .IN2(n1419), .QN(n1418) );
  IBUFFX16 U2099 ( .INP(n1585), .ZN(n2017) );
  AOI22X1 U2100 ( .IN1(n1944), .IN2(n2107), .IN3(n2087), .IN4(n1943), .QN(
        n1899) );
  INVX0 U2101 ( .INP(n1594), .ZN(n1900) );
  INVX0 U2102 ( .INP(n1900), .ZN(n1901) );
  OA22X1 U2103 ( .IN1(n1601), .IN2(n1057), .IN3(n2018), .IN4(n1174), .Q(n1600)
         );
  INVX0 U2104 ( .INP(g638), .ZN(n1902) );
  NAND3X1 U2105 ( .IN1(n1137), .IN2(n1993), .IN3(n1485), .QN(n1290) );
  NBUFFX2 U2106 ( .INP(n1587), .Z(n1919) );
  NBUFFX2 U2107 ( .INP(n1539), .Z(n1904) );
  AO21X1 U2108 ( .IN1(g594), .IN2(n1545), .IN3(n1249), .Q(n1906) );
  NAND2X0 U2109 ( .IN1(n2032), .IN2(n2031), .QN(n1907) );
  NAND2X0 U2110 ( .IN1(n2032), .IN2(n2031), .QN(n2041) );
  OR2X1 U2111 ( .IN1(n1207), .IN2(g128), .Q(n1689) );
  INVX0 U2112 ( .INP(n2054), .ZN(n1908) );
  INVX0 U2113 ( .INP(n1617), .ZN(n1917) );
  NBUFFX2 U2114 ( .INP(g694), .Z(n1909) );
  NBUFFX2 U2115 ( .INP(n1200), .Z(n1910) );
  NBUFFX2 U2116 ( .INP(n1200), .Z(n1911) );
  NBUFFX2 U2117 ( .INP(n1679), .Z(n1913) );
  INVX0 U2118 ( .INP(n1865), .ZN(n1965) );
  NBUFFX2 U2119 ( .INP(n1793), .Z(n2100) );
  INVX0 U2120 ( .INP(n1947), .ZN(n1618) );
  OA222X1 U2121 ( .IN1(n1895), .IN2(n1178), .IN3(n1809), .IN4(n1806), .IN5(
        n1168), .IN6(n1841), .Q(n1451) );
  NBUFFX2 U2122 ( .INP(g683), .Z(n1916) );
  NBUFFX2 U2123 ( .INP(g696), .Z(n1918) );
  AND2X1 U2124 ( .IN1(n1451), .IN2(n1450), .Q(n1921) );
  DELLN2X2 U2125 ( .INP(g28), .Z(n1923) );
  INVX0 U2126 ( .INP(n1590), .ZN(n1926) );
  INVX0 U2127 ( .INP(n1926), .ZN(n1927) );
  AOI22X1 U2128 ( .IN1(n2021), .IN2(n1894), .IN3(n1292), .IN4(n2044), .QN(
        n1264) );
  DELLN1X2 U2129 ( .INP(g658), .Z(n2044) );
  INVX0 U2130 ( .INP(n1129), .ZN(n1929) );
  OA21X1 U2131 ( .IN1(n1784), .IN2(n1569), .IN3(g676), .Q(n1483) );
  NAND3X1 U2132 ( .IN1(n1251), .IN2(n1252), .IN3(n1250), .QN(n1276) );
  INVX0 U2133 ( .INP(g685), .ZN(n1137) );
  NAND3X0 U2134 ( .IN1(n1453), .IN2(n1921), .IN3(n1452), .QN(g6481) );
  XNOR2X2 U2135 ( .IN1(g338), .IN2(n2078), .Q(n1658) );
  NOR4X1 U2136 ( .IN1(n1164), .IN2(g338), .IN3(g341), .IN4(g345), .QN(n1663)
         );
  DELLN2X2 U2137 ( .INP(n1569), .Z(n1930) );
  AND2X1 U2138 ( .IN1(n1374), .IN2(n1373), .Q(n1982) );
  AO21X1 U2139 ( .IN1(n1917), .IN2(n1612), .IN3(n1582), .Q(g6108) );
  AO21X1 U2140 ( .IN1(n1917), .IN2(n1596), .IN3(n1582), .Q(g6114) );
  AO21X1 U2141 ( .IN1(n1917), .IN2(n1606), .IN3(n1582), .Q(g6109) );
  INVX0 U2142 ( .INP(n1965), .ZN(n1931) );
  INVX0 U2143 ( .INP(n1965), .ZN(n1966) );
  XNOR2X1 U2144 ( .IN1(n1933), .IN2(n1128), .Q(n1636) );
  INVX0 U2145 ( .INP(n1091), .ZN(n1933) );
  INVX0 U2146 ( .INP(g278), .ZN(n1091) );
  AO21X1 U2147 ( .IN1(n1290), .IN2(n1482), .IN3(n1966), .Q(n1934) );
  AO22X1 U2148 ( .IN1(n1081), .IN2(n1952), .IN3(n1563), .IN4(n1885), .Q(g6289)
         );
  NAND4X0 U2149 ( .IN1(n1481), .IN2(n1167), .IN3(n1993), .IN4(n1086), .QN(
        n1935) );
  INVX0 U2150 ( .INP(g341), .ZN(n1936) );
  AND3X1 U2151 ( .IN1(n1460), .IN2(n1458), .IN3(n1449), .Q(n1937) );
  AND2X1 U2152 ( .IN1(n1472), .IN2(n1937), .Q(n1467) );
  AND3X1 U2153 ( .IN1(n1487), .IN2(n1938), .IN3(n1784), .Q(n1479) );
  INVX0 U2154 ( .INP(g204), .ZN(n1939) );
  NAND2X1 U2155 ( .IN1(n2027), .IN2(n1976), .QN(n1368) );
  NAND2X0 U2156 ( .IN1(n1392), .IN2(n1396), .QN(n1941) );
  NAND2X0 U2157 ( .IN1(n1392), .IN2(n1396), .QN(n1317) );
  AO22X1 U2158 ( .IN1(g465), .IN2(n1885), .IN3(n1081), .IN4(n1949), .Q(g6297)
         );
  AND2X1 U2159 ( .IN1(n1267), .IN2(n2023), .Q(n1942) );
  AND3X1 U2160 ( .IN1(n1982), .IN2(n1469), .IN3(n1935), .Q(n2027) );
  INVX0 U2161 ( .INP(n1414), .ZN(n1996) );
  OA221X1 U2162 ( .IN1(n1897), .IN2(n1173), .IN3(g489), .IN4(n1458), .IN5(
        n1459), .Q(n1457) );
  OA221X1 U2163 ( .IN1(n1897), .IN2(n1204), .IN3(g486), .IN4(n1458), .IN5(
        n1466), .Q(n1465) );
  XOR2X2 U2164 ( .IN1(n1139), .IN2(n2003), .Q(n1273) );
  NBUFFX2 U2165 ( .INP(n1468), .Z(n1946) );
  AND2X1 U2166 ( .IN1(n1133), .IN2(n1735), .Q(n1947) );
  NBUFFX2 U2167 ( .INP(n2044), .Z(n1948) );
  NAND2X1 U2168 ( .IN1(n1361), .IN2(n1362), .QN(n1349) );
  NBUFFX2 U2169 ( .INP(g691), .Z(n1949) );
  NBUFFX2 U2170 ( .INP(g682), .Z(n1950) );
  AO21X1 U2171 ( .IN1(n1588), .IN2(n1055), .IN3(n1893), .Q(g6116) );
  AO21X1 U2172 ( .IN1(n1581), .IN2(n1055), .IN3(n1893), .Q(g6118) );
  AO21X1 U2173 ( .IN1(n1599), .IN2(n1055), .IN3(n1893), .Q(g6113) );
  OA22X1 U2174 ( .IN1(g578), .IN2(n1149), .IN3(n1221), .IN4(n1196), .Q(n1578)
         );
  NBUFFX2 U2175 ( .INP(g693), .Z(n1952) );
  INVX0 U2176 ( .INP(n1953), .ZN(n1954) );
  XOR2X2 U2177 ( .IN1(n1403), .IN2(g478), .Q(n1386) );
  NAND3X0 U2178 ( .IN1(n1955), .IN2(n1956), .IN3(n1898), .QN(n1255) );
  OA22X1 U2179 ( .IN1(g161), .IN2(n1901), .IN3(n1855), .IN4(n1223), .Q(n1598)
         );
  AND2X1 U2180 ( .IN1(n1555), .IN2(g582), .Q(n1958) );
  AND2X1 U2181 ( .IN1(n1958), .IN2(n1959), .Q(n1545) );
  AND2X1 U2182 ( .IN1(g590), .IN2(n1727), .Q(n1959) );
  AO22X1 U2183 ( .IN1(n1048), .IN2(n1283), .IN3(n1284), .IN4(n2086), .Q(n1282)
         );
  INVX0 U2184 ( .INP(n2112), .ZN(n1960) );
  INVX0 U2185 ( .INP(n2112), .ZN(n1961) );
  AND2X1 U2186 ( .IN1(n1316), .IN2(n1317), .Q(n1962) );
  NAND2X1 U2187 ( .IN1(n1285), .IN2(n1799), .QN(n1963) );
  NAND2X0 U2188 ( .IN1(n1283), .IN2(n1117), .QN(n1964) );
  NAND3X0 U2189 ( .IN1(n1964), .IN2(n1963), .IN3(g260), .QN(n1284) );
  NOR2X0 U2190 ( .IN1(n2046), .IN2(n1742), .QN(g6291) );
  NAND2X1 U2191 ( .IN1(n1323), .IN2(n1744), .QN(n1322) );
  NAND2X0 U2192 ( .IN1(n1549), .IN2(n1727), .QN(n1546) );
  NBUFFX2 U2193 ( .INP(n1488), .Z(n1967) );
  NBUFFX2 U2194 ( .INP(n1475), .Z(n1969) );
  NBUFFX2 U2195 ( .INP(n1622), .Z(n1970) );
  NOR2X0 U2196 ( .IN1(n1666), .IN2(n1731), .QN(n1660) );
  NAND2X0 U2197 ( .IN1(n1467), .IN2(n1946), .QN(n1971) );
  INVX0 U2198 ( .INP(n1470), .ZN(n1972) );
  INVX0 U2199 ( .INP(n1470), .ZN(n1973) );
  NBUFFX2 U2200 ( .INP(n1431), .Z(n1974) );
  AND4X1 U2201 ( .IN1(n1472), .IN2(n1460), .IN3(n1449), .IN4(n1458), .Q(n1976)
         );
  AND3X1 U2202 ( .IN1(n1702), .IN2(n1701), .IN3(n1864), .Q(n1125) );
  AO21X1 U2203 ( .IN1(n1558), .IN2(n1559), .IN3(n1383), .Q(n1557) );
  INVX0 U2204 ( .INP(n1754), .ZN(n1979) );
  AOI22X1 U2205 ( .IN1(n1587), .IN2(n1118), .IN3(g188), .IN4(n1586), .QN(n1983) );
  AND2X1 U2206 ( .IN1(n2065), .IN2(g98), .Q(n1984) );
  AND2X1 U2207 ( .IN1(n1251), .IN2(n1984), .Q(n1271) );
  NAND2X0 U2208 ( .IN1(n1838), .IN2(n1853), .QN(n1393) );
  INVX0 U2209 ( .INP(n1949), .ZN(n1987) );
  AND3X1 U2210 ( .IN1(n1223), .IN2(n1112), .IN3(n1188), .Q(n1990) );
  XOR2X2 U2211 ( .IN1(n1821), .IN2(n1743), .Q(n1323) );
  XNOR2X1 U2212 ( .IN1(n1195), .IN2(n1991), .Q(n1497) );
  XOR2X1 U2213 ( .IN1(n1715), .IN2(g613), .Q(n1714) );
  NAND2X0 U2214 ( .IN1(n1594), .IN2(n1990), .QN(n1587) );
  INVX0 U2215 ( .INP(n1141), .ZN(n1992) );
  INVX0 U2216 ( .INP(n1994), .ZN(n1995) );
  INVX0 U2217 ( .INP(n1996), .ZN(n1997) );
  NOR2X0 U2218 ( .IN1(n1222), .IN2(n1129), .QN(n1414) );
  INVX0 U2219 ( .INP(n1381), .ZN(n1131) );
  NBUFFX2 U2220 ( .INP(n2051), .Z(n2110) );
  INVX0 U2221 ( .INP(n1256), .ZN(n1104) );
  INVX0 U2222 ( .INP(n2112), .ZN(n2113) );
  INVX0 U2223 ( .INP(n2112), .ZN(n2114) );
  NBUFFX2 U2224 ( .INP(n1347), .Z(n2101) );
  INVX0 U2225 ( .INP(n1553), .ZN(n1080) );
  INVX0 U2226 ( .INP(n2076), .ZN(n1109) );
  INVX0 U2227 ( .INP(n1513), .ZN(n1120) );
  NBUFFX2 U2228 ( .INP(n1206), .Z(n2106) );
  NBUFFX2 U2229 ( .INP(n1206), .Z(n2108) );
  NBUFFX2 U2230 ( .INP(n1490), .Z(n2099) );
  NBUFFX2 U2231 ( .INP(n1490), .Z(n2098) );
  INVX0 U2232 ( .INP(n1291), .ZN(n1159) );
  NBUFFX2 U2233 ( .INP(n1206), .Z(n2107) );
  INVX0 U2234 ( .INP(n2081), .ZN(n1135) );
  INVX0 U2235 ( .INP(n1106), .ZN(n2018) );
  INVX0 U2236 ( .INP(g1802), .ZN(n1233) );
  INVX0 U2237 ( .INP(n1653), .ZN(n1152) );
  AND3X1 U2238 ( .IN1(n1615), .IN2(n1614), .IN3(n1977), .Q(n2068) );
  INVX0 U2239 ( .INP(n1645), .ZN(n1105) );
  NOR2X0 U2240 ( .IN1(n1306), .IN2(n1718), .QN(g3454) );
  AOI21X1 U2241 ( .IN1(n1325), .IN2(n1244), .IN3(n1538), .QN(n1998) );
  AO21X1 U2242 ( .IN1(n1543), .IN2(n1090), .IN3(n2046), .Q(g6437) );
  NAND2X0 U2243 ( .IN1(n1426), .IN2(n1149), .QN(n1423) );
  NAND2X0 U2244 ( .IN1(n1410), .IN2(n1149), .QN(n1408) );
  INVX0 U2245 ( .INP(n1389), .ZN(n1097) );
  INVX0 U2246 ( .INP(n1162), .ZN(n2112) );
  INVX0 U2247 ( .INP(g6791), .ZN(n1066) );
  INVX0 U2248 ( .INP(g5533), .ZN(n1063) );
  INVX0 U2249 ( .INP(g6793), .ZN(n1073) );
  INVX0 U2250 ( .INP(g5535), .ZN(n1096) );
  INVX0 U2251 ( .INP(g5625), .ZN(n1095) );
  INVX0 U2252 ( .INP(g5626), .ZN(n1059) );
  INVX0 U2253 ( .INP(n1551), .ZN(n1081) );
  INVX0 U2254 ( .INP(g598), .ZN(n1110) );
  AO22X1 U2255 ( .IN1(n2088), .IN2(n1856), .IN3(n1080), .IN4(n2021), .Q(g6287)
         );
  OA22X1 U2256 ( .IN1(n1184), .IN2(n2086), .IN3(n1119), .IN4(n2110), .Q(n1283)
         );
  INVX0 U2257 ( .INP(n1615), .ZN(n1230) );
  INVX0 U2258 ( .INP(n2048), .ZN(n1248) );
  INVX0 U2259 ( .INP(n1443), .ZN(n1085) );
  INVX0 U2260 ( .INP(n1794), .ZN(n1206) );
  INVX0 U2261 ( .INP(n1356), .ZN(n1192) );
  INVX0 U2262 ( .INP(n1355), .ZN(n1108) );
  INVX0 U2263 ( .INP(g5629), .ZN(n1065) );
  INVX0 U2264 ( .INP(g5628), .ZN(n1092) );
  INVX0 U2265 ( .INP(n1436), .ZN(n1072) );
  NAND2X0 U2266 ( .IN1(n1381), .IN2(n1659), .QN(g5303) );
  INVX0 U2267 ( .INP(n1402), .ZN(n1146) );
  INVX0 U2268 ( .INP(n1473), .ZN(n1084) );
  INVX0 U2269 ( .INP(n1857), .ZN(n2050) );
  NBUFFX2 U2270 ( .INP(n1869), .Z(n2102) );
  NBUFFX2 U2271 ( .INP(n1869), .Z(n2103) );
  NAND2X1 U2272 ( .IN1(n2092), .IN2(n1432), .QN(g6110) );
  NAND2X1 U2273 ( .IN1(n2094), .IN2(n1158), .QN(g6189) );
  NAND2X1 U2274 ( .IN1(n2093), .IN2(n1166), .QN(g6185) );
  NAND2X1 U2275 ( .IN1(n2092), .IN2(n1116), .QN(g6173) );
  INVX0 U2276 ( .INP(n1430), .ZN(n1123) );
  NOR2X0 U2277 ( .IN1(n1242), .IN2(n1243), .QN(n1329) );
  INVX0 U2278 ( .INP(n1471), .ZN(n1050) );
  INVX0 U2279 ( .INP(n2047), .ZN(n2049) );
  NBUFFX2 U2280 ( .INP(n1570), .Z(n2094) );
  NBUFFX2 U2281 ( .INP(n1570), .Z(n2093) );
  NBUFFX2 U2282 ( .INP(n1570), .Z(n2092) );
  NOR2X0 U2283 ( .IN1(n1875), .IN2(n2066), .QN(g1802) );
  NAND2X1 U2284 ( .IN1(n1275), .IN2(n1261), .QN(n1274) );
  NOR2X0 U2285 ( .IN1(n1229), .IN2(n1226), .QN(n1511) );
  INVX0 U2286 ( .INP(n2042), .ZN(n2043) );
  INVX0 U2287 ( .INP(n2030), .ZN(n1121) );
  INVX0 U2288 ( .INP(n1253), .ZN(n1078) );
  NBUFFX2 U2289 ( .INP(g610), .Z(n2039) );
  INVX0 U2290 ( .INP(n1432), .ZN(n1115) );
  INVX0 U2291 ( .INP(g209), .ZN(n1194) );
  INVX0 U2292 ( .INP(g638), .ZN(n1190) );
  NAND2X0 U2293 ( .IN1(n1398), .IN2(n1123), .QN(n1397) );
  INVX0 U2294 ( .INP(g410), .ZN(n1156) );
  INVX0 U2295 ( .INP(g5627), .ZN(n1093) );
  INVX0 U2296 ( .INP(g5624), .ZN(n1062) );
  INVX0 U2297 ( .INP(g402), .ZN(n1154) );
  INVX0 U2298 ( .INP(g461), .ZN(n1077) );
  INVX0 U2299 ( .INP(g5532), .ZN(n1094) );
  AND3X1 U2300 ( .IN1(n1258), .IN2(n1058), .IN3(n1259), .Q(n1257) );
  INVX0 U2301 ( .INP(g449), .ZN(n1142) );
  INVX0 U2302 ( .INP(g301), .ZN(n1238) );
  NAND2X0 U2303 ( .IN1(g516), .IN2(n1085), .QN(n1438) );
  NAND2X0 U2304 ( .IN1(n1592), .IN2(n1593), .QN(n1591) );
  INVX0 U2305 ( .INP(g193), .ZN(n1214) );
  INVX0 U2306 ( .INP(g166), .ZN(n1174) );
  INVX0 U2307 ( .INP(g341), .ZN(n1181) );
  INVX0 U2308 ( .INP(g188), .ZN(n1118) );
  NBUFFX2 U2309 ( .INP(g269), .Z(n2089) );
  INVX0 U2310 ( .INP(g205), .ZN(n1205) );
  OA21X1 U2311 ( .IN1(n1638), .IN2(n1639), .IN3(n1064), .Q(n1637) );
  AO22X1 U2312 ( .IN1(g374), .IN2(n1980), .IN3(n1526), .IN4(n1859), .Q(n1525)
         );
  AO222X1 U2313 ( .IN1(n1120), .IN2(n1506), .IN3(n1507), .IN4(n1148), .IN5(
        g390), .IN6(n1981), .Q(n1505) );
  NOR3X0 U2314 ( .IN1(n1190), .IN2(n1676), .IN3(n1678), .QN(g5017) );
  INVX0 U2315 ( .INP(g102), .ZN(n2065) );
  NOR2X0 U2316 ( .IN1(n1306), .IN2(g642), .QN(n1713) );
  INVX0 U2317 ( .INP(n2082), .ZN(n1245) );
  INVX0 U2318 ( .INP(g692), .ZN(n1221) );
  NAND2X0 U2319 ( .IN1(n1928), .IN2(n1167), .QN(n1482) );
  NOR2X0 U2320 ( .IN1(n1629), .IN2(n2106), .QN(n1628) );
  NOR2X0 U2321 ( .IN1(n1631), .IN2(n1122), .QN(n1630) );
  INVX0 U2322 ( .INP(g697), .ZN(n1139) );
  AO22X1 U2323 ( .IN1(g532), .IN2(n1885), .IN3(n1081), .IN4(n2021), .Q(g6301)
         );
  NOR2X0 U2324 ( .IN1(n2077), .IN2(n1663), .QN(n1661) );
  NAND2X1 U2325 ( .IN1(n1663), .IN2(n2078), .QN(n1662) );
  INVX0 U2326 ( .INP(g281), .ZN(n1145) );
  NOR2X0 U2327 ( .IN1(n1710), .IN2(n1902), .QN(g4219) );
  NOR2X0 U2328 ( .IN1(n1675), .IN2(n1902), .QN(g5149) );
  INVX0 U2329 ( .INP(g680), .ZN(n1184) );
  INVX0 U2330 ( .INP(g135), .ZN(n1215) );
  NAND2X0 U2331 ( .IN1(n1175), .IN2(n1564), .QN(n1563) );
  NOR2X0 U2332 ( .IN1(n1677), .IN2(n1131), .QN(g5050) );
  XNOR2X1 U2333 ( .IN1(n1989), .IN2(g353), .Q(n1677) );
  INVX0 U2334 ( .INP(g532), .ZN(n1225) );
  INVX0 U2335 ( .INP(g512), .ZN(n1224) );
  INVX0 U2336 ( .INP(g504), .ZN(n1173) );
  NOR4X0 U2337 ( .IN1(n1352), .IN2(n1350), .IN3(n1351), .IN4(n1349), .QN(n1342) );
  DELLN1X2 U2338 ( .INP(n1784), .Z(g4110) );
  NOR3X0 U2339 ( .IN1(n1908), .IN2(n1549), .IN3(n1554), .QN(g6295) );
  NOR2X0 U2340 ( .IN1(n1571), .IN2(n1572), .QN(g6142) );
  NOR4X0 U2341 ( .IN1(n1580), .IN2(n1213), .IN3(g590), .IN4(n1196), .QN(n1571)
         );
  OR2X1 U2342 ( .IN1(n1999), .IN2(n2000), .Q(n1526) );
  INVX0 U2343 ( .INP(g59), .ZN(n1229) );
  NOR2X0 U2344 ( .IN1(g332), .IN2(n1382), .QN(n1380) );
  NAND2X0 U2345 ( .IN1(n1291), .IN2(n1150), .QN(n1379) );
  NAND2X0 U2346 ( .IN1(n1658), .IN2(n1381), .QN(g5323) );
  INVX0 U2347 ( .INP(g695), .ZN(n1076) );
  INVX0 U2348 ( .INP(g683), .ZN(n1179) );
  INVX0 U2349 ( .INP(g280), .ZN(n1193) );
  INVX0 U2350 ( .INP(g696), .ZN(n1177) );
  INVX0 U2351 ( .INP(g694), .ZN(n1227) );
  INVX0 U2352 ( .INP(g332), .ZN(n1054) );
  NAND2X0 U2353 ( .IN1(n1111), .IN2(n1415), .QN(g6702) );
  NOR4X0 U2354 ( .IN1(n1295), .IN2(n1296), .IN3(n1297), .IN4(n1298), .QN(n1294) );
  INVX0 U2355 ( .INP(g353), .ZN(n1180) );
  INVX0 U2356 ( .INP(g357), .ZN(n1172) );
  INVX0 U2357 ( .INP(g6690), .ZN(n1147) );
  INVX0 U2358 ( .INP(g6684), .ZN(n1198) );
  NBUFFX2 U2359 ( .INP(g684), .Z(n2030) );
  NAND2X1 U2360 ( .IN1(n2094), .IN2(n1210), .QN(g6170) );
  INVX0 U2361 ( .INP(g6688), .ZN(n1210) );
  NAND2X1 U2362 ( .IN1(n2094), .IN2(n1211), .QN(g6179) );
  INVX0 U2363 ( .INP(g6691), .ZN(n1211) );
  NAND2X1 U2364 ( .IN1(n2093), .IN2(n1130), .QN(g6167) );
  INVX0 U2365 ( .INP(g6686), .ZN(n1130) );
  INVX0 U2366 ( .INP(g679), .ZN(n1182) );
  NAND2X0 U2367 ( .IN1(n1291), .IN2(n1318), .QN(n1266) );
  NOR2X0 U2368 ( .IN1(n2043), .IN2(n1248), .QN(n1314) );
  OR2X1 U2369 ( .IN1(n2001), .IN2(n2002), .Q(n1311) );
  AND3X1 U2370 ( .IN1(n2043), .IN2(n1248), .IN3(n1951), .Q(n2002) );
  INVX0 U2371 ( .INP(g678), .ZN(n1051) );
  AO221X1 U2372 ( .IN1(g135), .IN2(n1685), .IN3(n1686), .IN4(n1102), .IN5(
        n1104), .Q(g4752) );
  INVX0 U2373 ( .INP(n1687), .ZN(n1102) );
  INVX0 U2374 ( .INP(g606), .ZN(n1117) );
  INVX0 U2375 ( .INP(g143), .ZN(n1185) );
  INVX0 U2376 ( .INP(g170), .ZN(n1188) );
  INVX0 U2377 ( .INP(g152), .ZN(n1220) );
  INVX0 U2378 ( .INP(g161), .ZN(n1223) );
  AO22X1 U2379 ( .IN1(n1260), .IN2(n1278), .IN3(n1261), .IN4(g123), .Q(n2003)
         );
  NAND2X1 U2380 ( .IN1(n1682), .IN2(n1256), .QN(g4773) );
  NBUFFX2 U2381 ( .INP(g269), .Z(n2091) );
  NBUFFX2 U2382 ( .INP(g269), .Z(n2090) );
  INVX0 U2383 ( .INP(g677), .ZN(n1212) );
  INVX0 U2384 ( .INP(g206), .ZN(n1140) );
  INVX0 U2385 ( .INP(g123), .ZN(n1058) );
  INVX0 U2386 ( .INP(g207), .ZN(n2034) );
  INVX0 U2387 ( .INP(g22), .ZN(n1235) );
  NOR3X0 U2388 ( .IN1(n2036), .IN2(n2037), .IN3(n1673), .QN(g5167) );
  INVX0 U2389 ( .INP(g107), .ZN(n1234) );
  NBUFFX2 U2390 ( .INP(g323), .Z(n2078) );
  NBUFFX2 U2391 ( .INP(g345), .Z(n2077) );
  NOR3X0 U2392 ( .IN1(n1249), .IN2(n1712), .IN3(n1716), .QN(g3768) );
  INVX0 U2393 ( .INP(g208), .ZN(n1122) );
  INVX0 U2394 ( .INP(g465), .ZN(n1087) );
  INVX0 U2395 ( .INP(g6685), .ZN(n1166) );
  INVX0 U2396 ( .INP(g6687), .ZN(n1158) );
  INVX0 U2397 ( .INP(g6689), .ZN(n1116) );
  INVX0 U2398 ( .INP(g541), .ZN(n1175) );
  INVX0 U2399 ( .INP(g646), .ZN(n1119) );
  INVX0 U2400 ( .INP(g79), .ZN(n1195) );
  INVX0 U2401 ( .INP(g179), .ZN(n1112) );
  INVX0 U2402 ( .INP(g84), .ZN(n1088) );
  INVX0 U2403 ( .INP(g681), .ZN(n1126) );
  INVX0 U2404 ( .INP(g536), .ZN(n1178) );
  INVX0 U2405 ( .INP(g687), .ZN(n1171) );
  INVX0 U2406 ( .INP(g590), .ZN(n1113) );
  INVX0 U2407 ( .INP(g586), .ZN(n1165) );
  NAND2X0 U2408 ( .IN1(n1765), .IN2(n2067), .QN(n1260) );
  NOR3X0 U2409 ( .IN1(n2036), .IN2(n1986), .IN3(n1695), .QN(g4460) );
  NOR3X0 U2410 ( .IN1(n2036), .IN2(n1696), .IN3(n1711), .QN(g4157) );
  AOI21X1 U2411 ( .IN1(n1986), .IN2(g625), .IN3(g628), .QN(n1680) );
  NOR2X0 U2412 ( .IN1(n1689), .IN2(g131), .QN(n1686) );
  NOR2X0 U2413 ( .IN1(n1690), .IN2(n2036), .QN(g4687) );
  INVX0 U2414 ( .INP(g582), .ZN(n1213) );
  INVX0 U2415 ( .INP(g337), .ZN(n1150) );
  INVX0 U2416 ( .INP(g686), .ZN(n1189) );
  OR2X1 U2417 ( .IN1(g672), .IN2(n2004), .Q(g5231) );
  NOR3X0 U2418 ( .IN1(g22), .IN2(n2082), .IN3(n1930), .QN(n2004) );
  INVX0 U2419 ( .INP(g496), .ZN(n1111) );
  NOR2X0 U2420 ( .IN1(g266), .IN2(n1763), .QN(g3910) );
  INVX0 U2421 ( .INP(g492), .ZN(n1187) );
  INVX0 U2422 ( .INP(g323), .ZN(n1136) );
  NBUFFX2 U2423 ( .INP(n1783), .Z(n2082) );
  INVX0 U2424 ( .INP(g297), .ZN(n1155) );
  INVX0 U2425 ( .INP(g293), .ZN(n1168) );
  INVX0 U2426 ( .INP(g157), .ZN(n1138) );
  INVX0 U2427 ( .INP(g602), .ZN(n1191) );
  INVX0 U2428 ( .INP(g500), .ZN(n1204) );
  INVX0 U2429 ( .INP(g349), .ZN(n1164) );
  INVX0 U2430 ( .INP(g382), .ZN(n1216) );
  INVX0 U2431 ( .INP(g111), .ZN(n1209) );
  INVX0 U2432 ( .INP(g437), .ZN(n1127) );
  INVX0 U2433 ( .INP(g441), .ZN(n1163) );
  INVX0 U2434 ( .INP(g445), .ZN(n1170) );
  INVX0 U2435 ( .INP(g266), .ZN(n1219) );
  INVX0 U2436 ( .INP(g508), .ZN(n1202) );
  INVX0 U2437 ( .INP(g430), .ZN(n1157) );
  INVX0 U2438 ( .INP(g426), .ZN(n1143) );
  INVX0 U2439 ( .INP(g422), .ZN(n1197) );
  INVX0 U2440 ( .INP(g418), .ZN(n1153) );
  INVX0 U2441 ( .INP(g434), .ZN(n1218) );
  INVX0 U2442 ( .INP(g406), .ZN(n1203) );
  INVX0 U2443 ( .INP(g453), .ZN(n1161) );
  INVX0 U2444 ( .INP(g414), .ZN(n1217) );
  INVX0 U2445 ( .INP(g457), .ZN(n1151) );
  INVX0 U2446 ( .INP(g47), .ZN(n1247) );
  AO22X1 U2447 ( .IN1(n1949), .IN2(n1961), .IN3(n1640), .IN4(n1635), .Q(g5625)
         );
  NBUFFX2 U2448 ( .INP(g5468), .Z(g4307) );
  NBUFFX2 U2449 ( .INP(g5469), .Z(g4321) );
  NBUFFX2 U2450 ( .INP(g5137), .Z(g3600) );
  NBUFFX2 U2451 ( .INP(g705), .Z(g3222) );
  DELLN1X2 U2452 ( .INP(g564), .Z(g4422) );
  DELLN1X2 U2453 ( .INP(g47), .Z(g4112) );
  NBUFFX2 U2454 ( .INP(g44), .Z(g4107) );
  NBUFFX2 U2455 ( .INP(g23), .Z(g4098) );
  DELLN1X2 U2456 ( .INP(g22), .Z(g4104) );
  INVX0 U2457 ( .INP(n1639), .ZN(n1069) );
  NOR2X0 U2458 ( .IN1(n1160), .IN2(n1911), .QN(n1291) );
  INVX0 U2459 ( .INP(g691), .ZN(n1228) );
  AO221X1 U2460 ( .IN1(g693), .IN2(n1309), .IN3(n1310), .IN4(n2021), .IN5(
        n1311), .Q(n1308) );
  INVX0 U2461 ( .INP(g693), .ZN(n1149) );
  INVX0 U2462 ( .INP(n1079), .ZN(n2014) );
  INVX0 U2463 ( .INP(n2014), .ZN(n2015) );
  NOR2X0 U2464 ( .IN1(n1866), .IN2(n1236), .QN(n1381) );
  OA21X1 U2465 ( .IN1(n1633), .IN2(n1623), .IN3(n1889), .Q(n1632) );
  INVX0 U2466 ( .INP(n1538), .ZN(n1133) );
  INVX0 U2467 ( .INP(g277), .ZN(n1222) );
  INVX0 U2468 ( .INP(g690), .ZN(n2019) );
  INVX0 U2469 ( .INP(n2019), .ZN(n2020) );
  INVX0 U2470 ( .INP(n2019), .ZN(n2021) );
  INVX0 U2471 ( .INP(n1231), .ZN(n2022) );
  INVX0 U2472 ( .INP(n1254), .ZN(n1231) );
  INVX0 U2473 ( .INP(g338), .ZN(n1176) );
  NAND2X0 U2474 ( .IN1(n2093), .IN2(n1147), .QN(g6176) );
  NAND2X0 U2475 ( .IN1(n1187), .IN2(n1400), .QN(g6704) );
  OA21X1 U2476 ( .IN1(n1460), .IN2(n1187), .IN3(n1368), .Q(n1459) );
  OA21X1 U2477 ( .IN1(n1460), .IN2(n1111), .IN3(n1368), .Q(n1466) );
  NBUFFX2 U2478 ( .INP(n1236), .Z(n2026) );
  AO22X1 U2479 ( .IN1(n2016), .IN2(n1918), .IN3(g524), .IN4(n2097), .Q(g6310)
         );
  INVX0 U2480 ( .INP(n1567), .ZN(n1082) );
  NOR2X0 U2481 ( .IN1(n1179), .IN2(n1567), .QN(n1568) );
  NOR2X0 U2482 ( .IN1(g123), .IN2(n1876), .QN(n1278) );
  NBUFFX2 U2483 ( .INP(n2116), .Z(g1293) );
  NAND2X1 U2484 ( .IN1(n1714), .IN2(g639), .QN(g3828) );
  INVX0 U2485 ( .INP(g94), .ZN(n1251) );
  INVX0 U2486 ( .INP(g98), .ZN(n1252) );
  NOR2X0 U2487 ( .IN1(n1689), .IN2(g131), .QN(n2031) );
  AND2X1 U2488 ( .IN1(n2033), .IN2(n1215), .Q(n2032) );
  INVX0 U2489 ( .INP(g139), .ZN(n2033) );
  INVX0 U2490 ( .INP(g89), .ZN(n1250) );
  INVX0 U2491 ( .INP(n1442), .ZN(n1083) );
  OA221X1 U2492 ( .IN1(n1169), .IN2(n1442), .IN3(n1789), .IN4(n1932), .IN5(
        n1478), .Q(n1463) );
  OR2X1 U2493 ( .IN1(n2034), .IN2(n1194), .Q(n2035) );
  INVX0 U2494 ( .INP(g639), .ZN(n2036) );
  INVX0 U2495 ( .INP(g639), .ZN(n1249) );
  NBUFFX2 U2496 ( .INP(n1794), .Z(n2087) );
  NBUFFX2 U2497 ( .INP(g197), .Z(n2088) );
  NOR2X0 U2498 ( .IN1(n1293), .IN2(n1294), .QN(n1292) );
  OA21X1 U2499 ( .IN1(n1141), .IN2(g207), .IN3(n1631), .Q(n1638) );
  NBUFFX2 U2500 ( .INP(n1562), .Z(n2037) );
  AND2X1 U2501 ( .IN1(g602), .IN2(g613), .Q(n2038) );
  AND2X1 U2502 ( .IN1(g610), .IN2(n2038), .Q(n1717) );
  INVX0 U2503 ( .INP(n1191), .ZN(n2040) );
  INVX0 U2504 ( .INP(g276), .ZN(n1129) );
  NOR2X0 U2505 ( .IN1(n1922), .IN2(n1929), .QN(n1410) );
  NOR2X0 U2506 ( .IN1(n1146), .IN2(n1100), .QN(n1651) );
  INVX0 U2507 ( .INP(n1950), .ZN(n1114) );
  NOR2X0 U2508 ( .IN1(g682), .IN2(g681), .QN(n1476) );
  NOR2X0 U2509 ( .IN1(n1394), .IN2(n1818), .QN(n1391) );
  AND2X1 U2510 ( .IN1(g698), .IN2(g689), .Q(n1485) );
  INVX0 U2511 ( .INP(g698), .ZN(n1167) );
  INVX0 U2512 ( .INP(n1928), .ZN(n1086) );
  INVX0 U2513 ( .INP(g598), .ZN(n2042) );
  NBUFFX2 U2514 ( .INP(n1550), .Z(n2095) );
  INVX0 U2515 ( .INP(n2095), .ZN(n1079) );
  AO22X1 U2516 ( .IN1(n2015), .IN2(n1810), .IN3(g520), .IN4(n2096), .Q(g6309)
         );
  AO22X1 U2517 ( .IN1(n2015), .IN2(n1944), .IN3(g528), .IN4(n2096), .Q(g6286)
         );
  NOR2X0 U2518 ( .IN1(n2037), .IN2(n1886), .QN(n1561) );
  NOR2X0 U2519 ( .IN1(n1939), .IN2(n1205), .QN(n1425) );
  NAND2X0 U2520 ( .IN1(n1207), .IN2(n1694), .QN(g4497) );
  NAND2X0 U2521 ( .IN1(g586), .IN2(n1549), .QN(n1548) );
  INVX0 U2522 ( .INP(n1395), .ZN(n1070) );
  OA21X1 U2523 ( .IN1(n1996), .IN2(n2020), .IN3(g278), .Q(n1409) );
  INVX0 U2524 ( .INP(n2020), .ZN(n1169) );
  NOR2X0 U2525 ( .IN1(g74), .IN2(g69), .QN(n1542) );
  NAND2X0 U2526 ( .IN1(n1286), .IN2(g606), .QN(n1285) );
  NAND2X0 U2527 ( .IN1(g679), .IN2(n1286), .QN(n1287) );
  AO22X1 U2528 ( .IN1(g678), .IN2(n1910), .IN3(g642), .IN4(n2086), .Q(n1286)
         );
  NOR2X0 U2529 ( .IN1(n1555), .IN2(g582), .QN(n1554) );
  AND2X1 U2530 ( .IN1(g631), .IN2(n1674), .Q(n1562) );
  NOR2X0 U2531 ( .IN1(g687), .IN2(n1865), .QN(n1481) );
  NBUFFX2 U2532 ( .INP(n1906), .Z(n2046) );
  INVX0 U2533 ( .INP(n2084), .ZN(n2051) );
  NAND2X0 U2534 ( .IN1(g131), .IN2(n1689), .QN(n1688) );
  INVX0 U2535 ( .INP(n1686), .ZN(n1103) );
  NAND2X0 U2536 ( .IN1(n1687), .IN2(n1871), .QN(n1685) );
  NAND2X0 U2537 ( .IN1(n1686), .IN2(n1215), .QN(n1684) );
  INVX0 U2538 ( .INP(g114), .ZN(n1207) );
  NAND2X0 U2539 ( .IN1(n1845), .IN2(n1957), .QN(n1626) );
  NOR2X0 U2540 ( .IN1(n1957), .IN2(n1634), .QN(n1633) );
  OR2X1 U2541 ( .IN1(n1241), .IN2(n1842), .Q(n1326) );
  INVX0 U2542 ( .INP(n1590), .ZN(n1057) );
  INVX0 U2543 ( .INP(g567), .ZN(n2047) );
  INVX0 U2544 ( .INP(n2047), .ZN(n2048) );
  OA21X1 U2545 ( .IN1(n1117), .IN2(n2076), .IN3(n1119), .Q(n1692) );
  NOR2X0 U2546 ( .IN1(n1683), .IN2(n1902), .QN(g4761) );
  INVX0 U2547 ( .INP(g314), .ZN(n2069) );
  NAND2X0 U2548 ( .IN1(n1547), .IN2(n2054), .QN(g6426) );
  NAND2X0 U2549 ( .IN1(n2092), .IN2(n1198), .QN(g6182) );
  NAND2X0 U2550 ( .IN1(n1496), .IN2(n1844), .QN(n1493) );
  NOR2X0 U2551 ( .IN1(n1819), .IN2(g631), .QN(n1673) );
  NOR2X0 U2552 ( .IN1(n1712), .IN2(g619), .QN(n1711) );
  INVX0 U2553 ( .INP(n2115), .ZN(n2055) );
  INVX0 U2554 ( .INP(n2055), .ZN(n2057) );
  INVX0 U2555 ( .INP(n2056), .ZN(n2058) );
  INVX0 U2556 ( .INP(n2056), .ZN(n2059) );
  INVX0 U2557 ( .INP(n2056), .ZN(n2060) );
  INVX0 U2558 ( .INP(n1873), .ZN(n2061) );
  INVX0 U2559 ( .INP(n1873), .ZN(n2062) );
  INVX0 U2560 ( .INP(n2115), .ZN(n2063) );
  INVX0 U2561 ( .INP(n1697), .ZN(n1124) );
  NAND2X0 U2562 ( .IN1(g520), .IN2(n1085), .QN(n1433) );
  NOR2X0 U2563 ( .IN1(n1978), .IN2(n2050), .QN(n1722) );
  NAND2X0 U2564 ( .IN1(n1136), .IN2(n1691), .QN(g4607) );
  NOR2X0 U2565 ( .IN1(n2026), .IN2(n1240), .QN(n1534) );
  INVX0 U2566 ( .INP(n1232), .ZN(n2066) );
  OA21X1 U2567 ( .IN1(g148), .IN2(n2018), .IN3(n1056), .Q(n1616) );
  NOR2X0 U2568 ( .IN1(n1607), .IN2(n2017), .QN(n1590) );
  NOR2X0 U2569 ( .IN1(n2017), .IN2(n1614), .QN(n1607) );
  NOR2X0 U2570 ( .IN1(n1997), .IN2(n1816), .QN(n1640) );
  NAND2X0 U2571 ( .IN1(n1390), .IN2(n1101), .QN(n1387) );
  AND2X1 U2572 ( .IN1(n1613), .IN2(n2068), .Q(n1582) );
  NOR2X0 U2573 ( .IN1(n1696), .IN2(g622), .QN(n1695) );
  OA21X1 U2574 ( .IN1(n1985), .IN2(g594), .IN3(n2054), .Q(g6304) );
  NOR2X0 U2575 ( .IN1(n2039), .IN2(n1191), .QN(n1719) );
  INVX0 U2576 ( .INP(n1985), .ZN(n1090) );
  INVX0 U2577 ( .INP(n1617), .ZN(n1055) );
  NAND3X1 U2578 ( .IN1(n1122), .IN2(n1087), .IN3(n1560), .QN(n1558) );
  NOR2X0 U2579 ( .IN1(n1896), .IN2(n1426), .QN(n1644) );
  OA21X1 U2580 ( .IN1(n1896), .IN2(g206), .IN3(n1992), .Q(n1641) );
  NAND2X0 U2581 ( .IN1(g208), .IN2(n1560), .QN(n1395) );
  NOR2X0 U2582 ( .IN1(n1430), .IN2(n1560), .QN(n1431) );
  NOR2X0 U2583 ( .IN1(n1872), .IN2(n1940), .QN(n1426) );
  NAND2X0 U2584 ( .IN1(g206), .IN2(n1425), .QN(n1643) );
  INVX0 U2585 ( .INP(n1752), .ZN(n1241) );
  NOR2X0 U2586 ( .IN1(n1762), .IN2(n2052), .QN(n1539) );
  INVX0 U2587 ( .INP(n1388), .ZN(n1101) );
  NOR2X0 U2588 ( .IN1(n1901), .IN2(n1855), .QN(n1601) );
  NAND2X0 U2589 ( .IN1(n1760), .IN2(n1232), .QN(n1261) );
  NOR2X0 U2590 ( .IN1(n1552), .IN2(n2046), .QN(g6299) );
  NOR2X0 U2591 ( .IN1(n1717), .IN2(g616), .QN(n1716) );
  NAND2X0 U2592 ( .IN1(n1113), .IN2(n1546), .QN(n1543) );
  NOR2X0 U2593 ( .IN1(n1249), .IN2(n2040), .QN(g2861) );
  NAND2X0 U2594 ( .IN1(n2039), .IN2(n2040), .QN(n1715) );
  INVX0 U2595 ( .INP(n1321), .ZN(n1236) );
  NAND2X0 U2596 ( .IN1(n1467), .IN2(n1468), .QN(n2072) );
  NAND2X0 U2597 ( .IN1(n1467), .IN2(n1946), .QN(n2073) );
  OA21X1 U2598 ( .IN1(g662), .IN2(g266), .IN3(n2051), .Q(n1487) );
  NOR2X0 U2599 ( .IN1(n2049), .IN2(g598), .QN(n1310) );
  NOR2X0 U2600 ( .IN1(n2049), .IN2(n1110), .QN(n1315) );
  NAND2X0 U2601 ( .IN1(g638), .IN2(n2049), .QN(g3599) );
  NOR2X0 U2602 ( .IN1(n1820), .IN2(n1259), .QN(n1256) );
  OA21X1 U2603 ( .IN1(n2022), .IN2(n1230), .IN3(n1617), .Q(n1619) );
  NOR2X0 U2604 ( .IN1(n2024), .IN2(n2066), .QN(n1254) );
  NOR2X0 U2605 ( .IN1(n1948), .IN2(n1763), .QN(g3814) );
  NBUFFX2 U2606 ( .INP(g658), .Z(n2084) );
  NAND2X0 U2607 ( .IN1(g642), .IN2(n1306), .QN(n1693) );
  NAND2X0 U2608 ( .IN1(g378), .IN2(n1979), .QN(n1520) );
  OA21X1 U2609 ( .IN1(g366), .IN2(n1859), .IN3(n1494), .Q(n1536) );
  NAND3X1 U2610 ( .IN1(g681), .IN2(n1114), .IN3(n1969), .QN(n1473) );
  INVX0 U2611 ( .INP(n2075), .ZN(n1240) );
  NAND2X0 U2612 ( .IN1(n2089), .IN2(n1625), .QN(n1624) );
  INVX0 U2613 ( .INP(n2089), .ZN(n1162) );
  INVX0 U2614 ( .INP(n1124), .ZN(n2115) );
  NAND2X0 U2615 ( .IN1(g524), .IN2(n1085), .QN(n1375) );
  INVX0 U2616 ( .INP(n1833), .ZN(n2080) );
  NAND2X0 U2617 ( .IN1(g528), .IN2(n1085), .QN(n1367) );
  NOR4X0 U2618 ( .IN1(n1703), .IN2(n1704), .IN3(n1706), .IN4(n1705), .QN(n1702) );
  IBUFFX16 U2619 ( .INP(n2342), .ZN(n2339) );
  IBUFFX16 U2620 ( .INP(n2339), .ZN(n2340) );
  IBUFFX16 U2621 ( .INP(n2339), .ZN(n2341) );
  DELLN2X2 U2622 ( .INP(test_se), .Z(n2342) );
endmodule

